`timescale 1ns/1ns
module sine_table_11x16
(input c,
 input      [10:0] angle,
 output reg [15:0] sine);

initial sine = 16'h0;

always @(posedge c) begin
  case (angle)
    11'd0: sine = 16'h0;
    11'd1: sine = 16'h64;
    11'd2: sine = 16'hc9;
    11'd3: sine = 16'h12d;
    11'd4: sine = 16'h192;
    11'd5: sine = 16'h1f6;
    11'd6: sine = 16'h25b;
    11'd7: sine = 16'h2bf;
    11'd8: sine = 16'h324;
    11'd9: sine = 16'h388;
    11'd10: sine = 16'h3ed;
    11'd11: sine = 16'h451;
    11'd12: sine = 16'h4b6;
    11'd13: sine = 16'h51a;
    11'd14: sine = 16'h57e;
    11'd15: sine = 16'h5e3;
    11'd16: sine = 16'h647;
    11'd17: sine = 16'h6ac;
    11'd18: sine = 16'h710;
    11'd19: sine = 16'h774;
    11'd20: sine = 16'h7d9;
    11'd21: sine = 16'h83d;
    11'd22: sine = 16'h8a1;
    11'd23: sine = 16'h906;
    11'd24: sine = 16'h96a;
    11'd25: sine = 16'h9ce;
    11'd26: sine = 16'ha32;
    11'd27: sine = 16'ha97;
    11'd28: sine = 16'hafb;
    11'd29: sine = 16'hb5f;
    11'd30: sine = 16'hbc3;
    11'd31: sine = 16'hc27;
    11'd32: sine = 16'hc8b;
    11'd33: sine = 16'hcef;
    11'd34: sine = 16'hd53;
    11'd35: sine = 16'hdb7;
    11'd36: sine = 16'he1b;
    11'd37: sine = 16'he7f;
    11'd38: sine = 16'hee3;
    11'd39: sine = 16'hf47;
    11'd40: sine = 16'hfab;
    11'd41: sine = 16'h100e;
    11'd42: sine = 16'h1072;
    11'd43: sine = 16'h10d6;
    11'd44: sine = 16'h1139;
    11'd45: sine = 16'h119d;
    11'd46: sine = 16'h1200;
    11'd47: sine = 16'h1264;
    11'd48: sine = 16'h12c7;
    11'd49: sine = 16'h132b;
    11'd50: sine = 16'h138e;
    11'd51: sine = 16'h13f2;
    11'd52: sine = 16'h1455;
    11'd53: sine = 16'h14b8;
    11'd54: sine = 16'h151b;
    11'd55: sine = 16'h157e;
    11'd56: sine = 16'h15e1;
    11'd57: sine = 16'h1644;
    11'd58: sine = 16'h16a7;
    11'd59: sine = 16'h170a;
    11'd60: sine = 16'h176d;
    11'd61: sine = 16'h17d0;
    11'd62: sine = 16'h1833;
    11'd63: sine = 16'h1895;
    11'd64: sine = 16'h18f8;
    11'd65: sine = 16'h195b;
    11'd66: sine = 16'h19bd;
    11'd67: sine = 16'h1a20;
    11'd68: sine = 16'h1a82;
    11'd69: sine = 16'h1ae4;
    11'd70: sine = 16'h1b46;
    11'd71: sine = 16'h1ba9;
    11'd72: sine = 16'h1c0b;
    11'd73: sine = 16'h1c6d;
    11'd74: sine = 16'h1ccf;
    11'd75: sine = 16'h1d31;
    11'd76: sine = 16'h1d93;
    11'd77: sine = 16'h1df4;
    11'd78: sine = 16'h1e56;
    11'd79: sine = 16'h1eb8;
    11'd80: sine = 16'h1f19;
    11'd81: sine = 16'h1f7b;
    11'd82: sine = 16'h1fdc;
    11'd83: sine = 16'h203d;
    11'd84: sine = 16'h209f;
    11'd85: sine = 16'h2100;
    11'd86: sine = 16'h2161;
    11'd87: sine = 16'h21c2;
    11'd88: sine = 16'h2223;
    11'd89: sine = 16'h2284;
    11'd90: sine = 16'h22e4;
    11'd91: sine = 16'h2345;
    11'd92: sine = 16'h23a6;
    11'd93: sine = 16'h2406;
    11'd94: sine = 16'h2467;
    11'd95: sine = 16'h24c7;
    11'd96: sine = 16'h2527;
    11'd97: sine = 16'h2587;
    11'd98: sine = 16'h25e7;
    11'd99: sine = 16'h2647;
    11'd100: sine = 16'h26a7;
    11'd101: sine = 16'h2707;
    11'd102: sine = 16'h2767;
    11'd103: sine = 16'h27c6;
    11'd104: sine = 16'h2826;
    11'd105: sine = 16'h2885;
    11'd106: sine = 16'h28e5;
    11'd107: sine = 16'h2944;
    11'd108: sine = 16'h29a3;
    11'd109: sine = 16'h2a02;
    11'd110: sine = 16'h2a61;
    11'd111: sine = 16'h2ac0;
    11'd112: sine = 16'h2b1e;
    11'd113: sine = 16'h2b7d;
    11'd114: sine = 16'h2bdb;
    11'd115: sine = 16'h2c3a;
    11'd116: sine = 16'h2c98;
    11'd117: sine = 16'h2cf6;
    11'd118: sine = 16'h2d54;
    11'd119: sine = 16'h2db2;
    11'd120: sine = 16'h2e10;
    11'd121: sine = 16'h2e6e;
    11'd122: sine = 16'h2ecc;
    11'd123: sine = 16'h2f29;
    11'd124: sine = 16'h2f86;
    11'd125: sine = 16'h2fe4;
    11'd126: sine = 16'h3041;
    11'd127: sine = 16'h309e;
    11'd128: sine = 16'h30fb;
    11'd129: sine = 16'h3158;
    11'd130: sine = 16'h31b4;
    11'd131: sine = 16'h3211;
    11'd132: sine = 16'h326d;
    11'd133: sine = 16'h32ca;
    11'd134: sine = 16'h3326;
    11'd135: sine = 16'h3382;
    11'd136: sine = 16'h33de;
    11'd137: sine = 16'h343a;
    11'd138: sine = 16'h3496;
    11'd139: sine = 16'h34f1;
    11'd140: sine = 16'h354d;
    11'd141: sine = 16'h35a8;
    11'd142: sine = 16'h3603;
    11'd143: sine = 16'h365e;
    11'd144: sine = 16'h36b9;
    11'd145: sine = 16'h3714;
    11'd146: sine = 16'h376f;
    11'd147: sine = 16'h37c9;
    11'd148: sine = 16'h3824;
    11'd149: sine = 16'h387e;
    11'd150: sine = 16'h38d8;
    11'd151: sine = 16'h3932;
    11'd152: sine = 16'h398c;
    11'd153: sine = 16'h39e6;
    11'd154: sine = 16'h3a3f;
    11'd155: sine = 16'h3a99;
    11'd156: sine = 16'h3af2;
    11'd157: sine = 16'h3b4b;
    11'd158: sine = 16'h3ba4;
    11'd159: sine = 16'h3bfd;
    11'd160: sine = 16'h3c56;
    11'd161: sine = 16'h3cae;
    11'd162: sine = 16'h3d07;
    11'd163: sine = 16'h3d5f;
    11'd164: sine = 16'h3db7;
    11'd165: sine = 16'h3e0f;
    11'd166: sine = 16'h3e67;
    11'd167: sine = 16'h3ebf;
    11'd168: sine = 16'h3f16;
    11'd169: sine = 16'h3f6e;
    11'd170: sine = 16'h3fc5;
    11'd171: sine = 16'h401c;
    11'd172: sine = 16'h4073;
    11'd173: sine = 16'h40ca;
    11'd174: sine = 16'h4120;
    11'd175: sine = 16'h4177;
    11'd176: sine = 16'h41cd;
    11'd177: sine = 16'h4223;
    11'd178: sine = 16'h4279;
    11'd179: sine = 16'h42cf;
    11'd180: sine = 16'h4325;
    11'd181: sine = 16'h437a;
    11'd182: sine = 16'h43d0;
    11'd183: sine = 16'h4425;
    11'd184: sine = 16'h447a;
    11'd185: sine = 16'h44cf;
    11'd186: sine = 16'h4523;
    11'd187: sine = 16'h4578;
    11'd188: sine = 16'h45cc;
    11'd189: sine = 16'h4620;
    11'd190: sine = 16'h4674;
    11'd191: sine = 16'h46c8;
    11'd192: sine = 16'h471c;
    11'd193: sine = 16'h476f;
    11'd194: sine = 16'h47c3;
    11'd195: sine = 16'h4816;
    11'd196: sine = 16'h4869;
    11'd197: sine = 16'h48bc;
    11'd198: sine = 16'h490e;
    11'd199: sine = 16'h4961;
    11'd200: sine = 16'h49b3;
    11'd201: sine = 16'h4a05;
    11'd202: sine = 16'h4a57;
    11'd203: sine = 16'h4aa9;
    11'd204: sine = 16'h4afa;
    11'd205: sine = 16'h4b4c;
    11'd206: sine = 16'h4b9d;
    11'd207: sine = 16'h4bee;
    11'd208: sine = 16'h4c3f;
    11'd209: sine = 16'h4c8f;
    11'd210: sine = 16'h4ce0;
    11'd211: sine = 16'h4d30;
    11'd212: sine = 16'h4d80;
    11'd213: sine = 16'h4dd0;
    11'd214: sine = 16'h4e20;
    11'd215: sine = 16'h4e6f;
    11'd216: sine = 16'h4ebf;
    11'd217: sine = 16'h4f0e;
    11'd218: sine = 16'h4f5d;
    11'd219: sine = 16'h4fac;
    11'd220: sine = 16'h4ffa;
    11'd221: sine = 16'h5049;
    11'd222: sine = 16'h5097;
    11'd223: sine = 16'h50e5;
    11'd224: sine = 16'h5133;
    11'd225: sine = 16'h5180;
    11'd226: sine = 16'h51ce;
    11'd227: sine = 16'h521b;
    11'd228: sine = 16'h5268;
    11'd229: sine = 16'h52b5;
    11'd230: sine = 16'h5301;
    11'd231: sine = 16'h534e;
    11'd232: sine = 16'h539a;
    11'd233: sine = 16'h53e6;
    11'd234: sine = 16'h5432;
    11'd235: sine = 16'h547d;
    11'd236: sine = 16'h54c9;
    11'd237: sine = 16'h5514;
    11'd238: sine = 16'h555f;
    11'd239: sine = 16'h55aa;
    11'd240: sine = 16'h55f4;
    11'd241: sine = 16'h563f;
    11'd242: sine = 16'h5689;
    11'd243: sine = 16'h56d3;
    11'd244: sine = 16'h571d;
    11'd245: sine = 16'h5766;
    11'd246: sine = 16'h57b0;
    11'd247: sine = 16'h57f9;
    11'd248: sine = 16'h5842;
    11'd249: sine = 16'h588a;
    11'd250: sine = 16'h58d3;
    11'd251: sine = 16'h591b;
    11'd252: sine = 16'h5963;
    11'd253: sine = 16'h59ab;
    11'd254: sine = 16'h59f3;
    11'd255: sine = 16'h5a3a;
    11'd256: sine = 16'h5a81;
    11'd257: sine = 16'h5ac8;
    11'd258: sine = 16'h5b0f;
    11'd259: sine = 16'h5b56;
    11'd260: sine = 16'h5b9c;
    11'd261: sine = 16'h5be2;
    11'd262: sine = 16'h5c28;
    11'd263: sine = 16'h5c6d;
    11'd264: sine = 16'h5cb3;
    11'd265: sine = 16'h5cf8;
    11'd266: sine = 16'h5d3d;
    11'd267: sine = 16'h5d82;
    11'd268: sine = 16'h5dc6;
    11'd269: sine = 16'h5e0b;
    11'd270: sine = 16'h5e4f;
    11'd271: sine = 16'h5e93;
    11'd272: sine = 16'h5ed6;
    11'd273: sine = 16'h5f1a;
    11'd274: sine = 16'h5f5d;
    11'd275: sine = 16'h5fa0;
    11'd276: sine = 16'h5fe2;
    11'd277: sine = 16'h6025;
    11'd278: sine = 16'h6067;
    11'd279: sine = 16'h60a9;
    11'd280: sine = 16'h60eb;
    11'd281: sine = 16'h612d;
    11'd282: sine = 16'h616e;
    11'd283: sine = 16'h61af;
    11'd284: sine = 16'h61f0;
    11'd285: sine = 16'h6230;
    11'd286: sine = 16'h6271;
    11'd287: sine = 16'h62b1;
    11'd288: sine = 16'h62f1;
    11'd289: sine = 16'h6330;
    11'd290: sine = 16'h6370;
    11'd291: sine = 16'h63af;
    11'd292: sine = 16'h63ee;
    11'd293: sine = 16'h642d;
    11'd294: sine = 16'h646b;
    11'd295: sine = 16'h64a9;
    11'd296: sine = 16'h64e7;
    11'd297: sine = 16'h6525;
    11'd298: sine = 16'h6562;
    11'd299: sine = 16'h65a0;
    11'd300: sine = 16'h65dd;
    11'd301: sine = 16'h6619;
    11'd302: sine = 16'h6656;
    11'd303: sine = 16'h6692;
    11'd304: sine = 16'h66ce;
    11'd305: sine = 16'h670a;
    11'd306: sine = 16'h6745;
    11'd307: sine = 16'h6781;
    11'd308: sine = 16'h67bc;
    11'd309: sine = 16'h67f7;
    11'd310: sine = 16'h6831;
    11'd311: sine = 16'h686b;
    11'd312: sine = 16'h68a5;
    11'd313: sine = 16'h68df;
    11'd314: sine = 16'h6919;
    11'd315: sine = 16'h6952;
    11'd316: sine = 16'h698b;
    11'd317: sine = 16'h69c4;
    11'd318: sine = 16'h69fc;
    11'd319: sine = 16'h6a34;
    11'd320: sine = 16'h6a6c;
    11'd321: sine = 16'h6aa4;
    11'd322: sine = 16'h6adb;
    11'd323: sine = 16'h6b13;
    11'd324: sine = 16'h6b4a;
    11'd325: sine = 16'h6b80;
    11'd326: sine = 16'h6bb7;
    11'd327: sine = 16'h6bed;
    11'd328: sine = 16'h6c23;
    11'd329: sine = 16'h6c58;
    11'd330: sine = 16'h6c8e;
    11'd331: sine = 16'h6cc3;
    11'd332: sine = 16'h6cf8;
    11'd333: sine = 16'h6d2c;
    11'd334: sine = 16'h6d61;
    11'd335: sine = 16'h6d95;
    11'd336: sine = 16'h6dc9;
    11'd337: sine = 16'h6dfc;
    11'd338: sine = 16'h6e30;
    11'd339: sine = 16'h6e63;
    11'd340: sine = 16'h6e95;
    11'd341: sine = 16'h6ec8;
    11'd342: sine = 16'h6efa;
    11'd343: sine = 16'h6f2c;
    11'd344: sine = 16'h6f5e;
    11'd345: sine = 16'h6f8f;
    11'd346: sine = 16'h6fc0;
    11'd347: sine = 16'h6ff1;
    11'd348: sine = 16'h7022;
    11'd349: sine = 16'h7052;
    11'd350: sine = 16'h7082;
    11'd351: sine = 16'h70b2;
    11'd352: sine = 16'h70e1;
    11'd353: sine = 16'h7111;
    11'd354: sine = 16'h7140;
    11'd355: sine = 16'h716e;
    11'd356: sine = 16'h719d;
    11'd357: sine = 16'h71cb;
    11'd358: sine = 16'h71f9;
    11'd359: sine = 16'h7226;
    11'd360: sine = 16'h7254;
    11'd361: sine = 16'h7281;
    11'd362: sine = 16'h72ae;
    11'd363: sine = 16'h72da;
    11'd364: sine = 16'h7306;
    11'd365: sine = 16'h7332;
    11'd366: sine = 16'h735e;
    11'd367: sine = 16'h7389;
    11'd368: sine = 16'h73b5;
    11'd369: sine = 16'h73df;
    11'd370: sine = 16'h740a;
    11'd371: sine = 16'h7434;
    11'd372: sine = 16'h745e;
    11'd373: sine = 16'h7488;
    11'd374: sine = 16'h74b1;
    11'd375: sine = 16'h74db;
    11'd376: sine = 16'h7503;
    11'd377: sine = 16'h752c;
    11'd378: sine = 16'h7554;
    11'd379: sine = 16'h757c;
    11'd380: sine = 16'h75a4;
    11'd381: sine = 16'h75cc;
    11'd382: sine = 16'h75f3;
    11'd383: sine = 16'h761a;
    11'd384: sine = 16'h7640;
    11'd385: sine = 16'h7667;
    11'd386: sine = 16'h768d;
    11'd387: sine = 16'h76b2;
    11'd388: sine = 16'h76d8;
    11'd389: sine = 16'h76fd;
    11'd390: sine = 16'h7722;
    11'd391: sine = 16'h7747;
    11'd392: sine = 16'h776b;
    11'd393: sine = 16'h778f;
    11'd394: sine = 16'h77b3;
    11'd395: sine = 16'h77d6;
    11'd396: sine = 16'h77f9;
    11'd397: sine = 16'h781c;
    11'd398: sine = 16'h783f;
    11'd399: sine = 16'h7861;
    11'd400: sine = 16'h7883;
    11'd401: sine = 16'h78a5;
    11'd402: sine = 16'h78c6;
    11'd403: sine = 16'h78e7;
    11'd404: sine = 16'h7908;
    11'd405: sine = 16'h7929;
    11'd406: sine = 16'h7949;
    11'd407: sine = 16'h7969;
    11'd408: sine = 16'h7989;
    11'd409: sine = 16'h79a8;
    11'd410: sine = 16'h79c7;
    11'd411: sine = 16'h79e6;
    11'd412: sine = 16'h7a04;
    11'd413: sine = 16'h7a23;
    11'd414: sine = 16'h7a41;
    11'd415: sine = 16'h7a5e;
    11'd416: sine = 16'h7a7c;
    11'd417: sine = 16'h7a99;
    11'd418: sine = 16'h7ab5;
    11'd419: sine = 16'h7ad2;
    11'd420: sine = 16'h7aee;
    11'd421: sine = 16'h7b0a;
    11'd422: sine = 16'h7b25;
    11'd423: sine = 16'h7b41;
    11'd424: sine = 16'h7b5c;
    11'd425: sine = 16'h7b76;
    11'd426: sine = 16'h7b91;
    11'd427: sine = 16'h7bab;
    11'd428: sine = 16'h7bc4;
    11'd429: sine = 16'h7bde;
    11'd430: sine = 16'h7bf7;
    11'd431: sine = 16'h7c10;
    11'd432: sine = 16'h7c29;
    11'd433: sine = 16'h7c41;
    11'd434: sine = 16'h7c59;
    11'd435: sine = 16'h7c70;
    11'd436: sine = 16'h7c88;
    11'd437: sine = 16'h7c9f;
    11'd438: sine = 16'h7cb6;
    11'd439: sine = 16'h7ccc;
    11'd440: sine = 16'h7ce2;
    11'd441: sine = 16'h7cf8;
    11'd442: sine = 16'h7d0e;
    11'd443: sine = 16'h7d23;
    11'd444: sine = 16'h7d38;
    11'd445: sine = 16'h7d4d;
    11'd446: sine = 16'h7d61;
    11'd447: sine = 16'h7d75;
    11'd448: sine = 16'h7d89;
    11'd449: sine = 16'h7d9c;
    11'd450: sine = 16'h7db0;
    11'd451: sine = 16'h7dc2;
    11'd452: sine = 16'h7dd5;
    11'd453: sine = 16'h7de7;
    11'd454: sine = 16'h7df9;
    11'd455: sine = 16'h7e0b;
    11'd456: sine = 16'h7e1c;
    11'd457: sine = 16'h7e2d;
    11'd458: sine = 16'h7e3e;
    11'd459: sine = 16'h7e4e;
    11'd460: sine = 16'h7e5e;
    11'd461: sine = 16'h7e6e;
    11'd462: sine = 16'h7e7e;
    11'd463: sine = 16'h7e8d;
    11'd464: sine = 16'h7e9c;
    11'd465: sine = 16'h7eaa;
    11'd466: sine = 16'h7eb9;
    11'd467: sine = 16'h7ec7;
    11'd468: sine = 16'h7ed4;
    11'd469: sine = 16'h7ee2;
    11'd470: sine = 16'h7eef;
    11'd471: sine = 16'h7efc;
    11'd472: sine = 16'h7f08;
    11'd473: sine = 16'h7f14;
    11'd474: sine = 16'h7f20;
    11'd475: sine = 16'h7f2c;
    11'd476: sine = 16'h7f37;
    11'd477: sine = 16'h7f42;
    11'd478: sine = 16'h7f4c;
    11'd479: sine = 16'h7f57;
    11'd480: sine = 16'h7f61;
    11'd481: sine = 16'h7f6a;
    11'd482: sine = 16'h7f74;
    11'd483: sine = 16'h7f7d;
    11'd484: sine = 16'h7f86;
    11'd485: sine = 16'h7f8e;
    11'd486: sine = 16'h7f96;
    11'd487: sine = 16'h7f9e;
    11'd488: sine = 16'h7fa6;
    11'd489: sine = 16'h7fad;
    11'd490: sine = 16'h7fb4;
    11'd491: sine = 16'h7fbb;
    11'd492: sine = 16'h7fc1;
    11'd493: sine = 16'h7fc7;
    11'd494: sine = 16'h7fcd;
    11'd495: sine = 16'h7fd2;
    11'd496: sine = 16'h7fd7;
    11'd497: sine = 16'h7fdc;
    11'd498: sine = 16'h7fe0;
    11'd499: sine = 16'h7fe4;
    11'd500: sine = 16'h7fe8;
    11'd501: sine = 16'h7fec;
    11'd502: sine = 16'h7fef;
    11'd503: sine = 16'h7ff2;
    11'd504: sine = 16'h7ff5;
    11'd505: sine = 16'h7ff7;
    11'd506: sine = 16'h7ff9;
    11'd507: sine = 16'h7ffb;
    11'd508: sine = 16'h7ffc;
    11'd509: sine = 16'h7ffd;
    11'd510: sine = 16'h7ffe;
    11'd511: sine = 16'h7ffe;
    11'd512: sine = 16'h7ffe;
    11'd513: sine = 16'h7ffe;
    11'd514: sine = 16'h7ffe;
    11'd515: sine = 16'h7ffd;
    11'd516: sine = 16'h7ffc;
    11'd517: sine = 16'h7ffb;
    11'd518: sine = 16'h7ff9;
    11'd519: sine = 16'h7ff7;
    11'd520: sine = 16'h7ff5;
    11'd521: sine = 16'h7ff2;
    11'd522: sine = 16'h7fef;
    11'd523: sine = 16'h7fec;
    11'd524: sine = 16'h7fe8;
    11'd525: sine = 16'h7fe4;
    11'd526: sine = 16'h7fe0;
    11'd527: sine = 16'h7fdc;
    11'd528: sine = 16'h7fd7;
    11'd529: sine = 16'h7fd2;
    11'd530: sine = 16'h7fcd;
    11'd531: sine = 16'h7fc7;
    11'd532: sine = 16'h7fc1;
    11'd533: sine = 16'h7fbb;
    11'd534: sine = 16'h7fb4;
    11'd535: sine = 16'h7fad;
    11'd536: sine = 16'h7fa6;
    11'd537: sine = 16'h7f9e;
    11'd538: sine = 16'h7f96;
    11'd539: sine = 16'h7f8e;
    11'd540: sine = 16'h7f86;
    11'd541: sine = 16'h7f7d;
    11'd542: sine = 16'h7f74;
    11'd543: sine = 16'h7f6a;
    11'd544: sine = 16'h7f61;
    11'd545: sine = 16'h7f57;
    11'd546: sine = 16'h7f4c;
    11'd547: sine = 16'h7f42;
    11'd548: sine = 16'h7f37;
    11'd549: sine = 16'h7f2c;
    11'd550: sine = 16'h7f20;
    11'd551: sine = 16'h7f14;
    11'd552: sine = 16'h7f08;
    11'd553: sine = 16'h7efc;
    11'd554: sine = 16'h7eef;
    11'd555: sine = 16'h7ee2;
    11'd556: sine = 16'h7ed4;
    11'd557: sine = 16'h7ec7;
    11'd558: sine = 16'h7eb9;
    11'd559: sine = 16'h7eaa;
    11'd560: sine = 16'h7e9c;
    11'd561: sine = 16'h7e8d;
    11'd562: sine = 16'h7e7e;
    11'd563: sine = 16'h7e6e;
    11'd564: sine = 16'h7e5e;
    11'd565: sine = 16'h7e4e;
    11'd566: sine = 16'h7e3e;
    11'd567: sine = 16'h7e2d;
    11'd568: sine = 16'h7e1c;
    11'd569: sine = 16'h7e0b;
    11'd570: sine = 16'h7df9;
    11'd571: sine = 16'h7de7;
    11'd572: sine = 16'h7dd5;
    11'd573: sine = 16'h7dc2;
    11'd574: sine = 16'h7db0;
    11'd575: sine = 16'h7d9c;
    11'd576: sine = 16'h7d89;
    11'd577: sine = 16'h7d75;
    11'd578: sine = 16'h7d61;
    11'd579: sine = 16'h7d4d;
    11'd580: sine = 16'h7d38;
    11'd581: sine = 16'h7d23;
    11'd582: sine = 16'h7d0e;
    11'd583: sine = 16'h7cf8;
    11'd584: sine = 16'h7ce2;
    11'd585: sine = 16'h7ccc;
    11'd586: sine = 16'h7cb6;
    11'd587: sine = 16'h7c9f;
    11'd588: sine = 16'h7c88;
    11'd589: sine = 16'h7c70;
    11'd590: sine = 16'h7c59;
    11'd591: sine = 16'h7c41;
    11'd592: sine = 16'h7c29;
    11'd593: sine = 16'h7c10;
    11'd594: sine = 16'h7bf7;
    11'd595: sine = 16'h7bde;
    11'd596: sine = 16'h7bc4;
    11'd597: sine = 16'h7bab;
    11'd598: sine = 16'h7b91;
    11'd599: sine = 16'h7b76;
    11'd600: sine = 16'h7b5c;
    11'd601: sine = 16'h7b41;
    11'd602: sine = 16'h7b25;
    11'd603: sine = 16'h7b0a;
    11'd604: sine = 16'h7aee;
    11'd605: sine = 16'h7ad2;
    11'd606: sine = 16'h7ab5;
    11'd607: sine = 16'h7a99;
    11'd608: sine = 16'h7a7c;
    11'd609: sine = 16'h7a5e;
    11'd610: sine = 16'h7a41;
    11'd611: sine = 16'h7a23;
    11'd612: sine = 16'h7a04;
    11'd613: sine = 16'h79e6;
    11'd614: sine = 16'h79c7;
    11'd615: sine = 16'h79a8;
    11'd616: sine = 16'h7989;
    11'd617: sine = 16'h7969;
    11'd618: sine = 16'h7949;
    11'd619: sine = 16'h7929;
    11'd620: sine = 16'h7908;
    11'd621: sine = 16'h78e7;
    11'd622: sine = 16'h78c6;
    11'd623: sine = 16'h78a5;
    11'd624: sine = 16'h7883;
    11'd625: sine = 16'h7861;
    11'd626: sine = 16'h783f;
    11'd627: sine = 16'h781c;
    11'd628: sine = 16'h77f9;
    11'd629: sine = 16'h77d6;
    11'd630: sine = 16'h77b3;
    11'd631: sine = 16'h778f;
    11'd632: sine = 16'h776b;
    11'd633: sine = 16'h7747;
    11'd634: sine = 16'h7722;
    11'd635: sine = 16'h76fd;
    11'd636: sine = 16'h76d8;
    11'd637: sine = 16'h76b2;
    11'd638: sine = 16'h768d;
    11'd639: sine = 16'h7667;
    11'd640: sine = 16'h7640;
    11'd641: sine = 16'h761a;
    11'd642: sine = 16'h75f3;
    11'd643: sine = 16'h75cc;
    11'd644: sine = 16'h75a4;
    11'd645: sine = 16'h757c;
    11'd646: sine = 16'h7554;
    11'd647: sine = 16'h752c;
    11'd648: sine = 16'h7503;
    11'd649: sine = 16'h74db;
    11'd650: sine = 16'h74b1;
    11'd651: sine = 16'h7488;
    11'd652: sine = 16'h745e;
    11'd653: sine = 16'h7434;
    11'd654: sine = 16'h740a;
    11'd655: sine = 16'h73df;
    11'd656: sine = 16'h73b5;
    11'd657: sine = 16'h7389;
    11'd658: sine = 16'h735e;
    11'd659: sine = 16'h7332;
    11'd660: sine = 16'h7306;
    11'd661: sine = 16'h72da;
    11'd662: sine = 16'h72ae;
    11'd663: sine = 16'h7281;
    11'd664: sine = 16'h7254;
    11'd665: sine = 16'h7226;
    11'd666: sine = 16'h71f9;
    11'd667: sine = 16'h71cb;
    11'd668: sine = 16'h719d;
    11'd669: sine = 16'h716e;
    11'd670: sine = 16'h7140;
    11'd671: sine = 16'h7111;
    11'd672: sine = 16'h70e1;
    11'd673: sine = 16'h70b2;
    11'd674: sine = 16'h7082;
    11'd675: sine = 16'h7052;
    11'd676: sine = 16'h7022;
    11'd677: sine = 16'h6ff1;
    11'd678: sine = 16'h6fc0;
    11'd679: sine = 16'h6f8f;
    11'd680: sine = 16'h6f5e;
    11'd681: sine = 16'h6f2c;
    11'd682: sine = 16'h6efa;
    11'd683: sine = 16'h6ec8;
    11'd684: sine = 16'h6e95;
    11'd685: sine = 16'h6e63;
    11'd686: sine = 16'h6e30;
    11'd687: sine = 16'h6dfc;
    11'd688: sine = 16'h6dc9;
    11'd689: sine = 16'h6d95;
    11'd690: sine = 16'h6d61;
    11'd691: sine = 16'h6d2c;
    11'd692: sine = 16'h6cf8;
    11'd693: sine = 16'h6cc3;
    11'd694: sine = 16'h6c8e;
    11'd695: sine = 16'h6c58;
    11'd696: sine = 16'h6c23;
    11'd697: sine = 16'h6bed;
    11'd698: sine = 16'h6bb7;
    11'd699: sine = 16'h6b80;
    11'd700: sine = 16'h6b4a;
    11'd701: sine = 16'h6b13;
    11'd702: sine = 16'h6adb;
    11'd703: sine = 16'h6aa4;
    11'd704: sine = 16'h6a6c;
    11'd705: sine = 16'h6a34;
    11'd706: sine = 16'h69fc;
    11'd707: sine = 16'h69c4;
    11'd708: sine = 16'h698b;
    11'd709: sine = 16'h6952;
    11'd710: sine = 16'h6919;
    11'd711: sine = 16'h68df;
    11'd712: sine = 16'h68a5;
    11'd713: sine = 16'h686b;
    11'd714: sine = 16'h6831;
    11'd715: sine = 16'h67f7;
    11'd716: sine = 16'h67bc;
    11'd717: sine = 16'h6781;
    11'd718: sine = 16'h6745;
    11'd719: sine = 16'h670a;
    11'd720: sine = 16'h66ce;
    11'd721: sine = 16'h6692;
    11'd722: sine = 16'h6656;
    11'd723: sine = 16'h6619;
    11'd724: sine = 16'h65dd;
    11'd725: sine = 16'h65a0;
    11'd726: sine = 16'h6562;
    11'd727: sine = 16'h6525;
    11'd728: sine = 16'h64e7;
    11'd729: sine = 16'h64a9;
    11'd730: sine = 16'h646b;
    11'd731: sine = 16'h642d;
    11'd732: sine = 16'h63ee;
    11'd733: sine = 16'h63af;
    11'd734: sine = 16'h6370;
    11'd735: sine = 16'h6330;
    11'd736: sine = 16'h62f1;
    11'd737: sine = 16'h62b1;
    11'd738: sine = 16'h6271;
    11'd739: sine = 16'h6230;
    11'd740: sine = 16'h61f0;
    11'd741: sine = 16'h61af;
    11'd742: sine = 16'h616e;
    11'd743: sine = 16'h612d;
    11'd744: sine = 16'h60eb;
    11'd745: sine = 16'h60a9;
    11'd746: sine = 16'h6067;
    11'd747: sine = 16'h6025;
    11'd748: sine = 16'h5fe2;
    11'd749: sine = 16'h5fa0;
    11'd750: sine = 16'h5f5d;
    11'd751: sine = 16'h5f1a;
    11'd752: sine = 16'h5ed6;
    11'd753: sine = 16'h5e93;
    11'd754: sine = 16'h5e4f;
    11'd755: sine = 16'h5e0b;
    11'd756: sine = 16'h5dc6;
    11'd757: sine = 16'h5d82;
    11'd758: sine = 16'h5d3d;
    11'd759: sine = 16'h5cf8;
    11'd760: sine = 16'h5cb3;
    11'd761: sine = 16'h5c6d;
    11'd762: sine = 16'h5c28;
    11'd763: sine = 16'h5be2;
    11'd764: sine = 16'h5b9c;
    11'd765: sine = 16'h5b56;
    11'd766: sine = 16'h5b0f;
    11'd767: sine = 16'h5ac8;
    11'd768: sine = 16'h5a81;
    11'd769: sine = 16'h5a3a;
    11'd770: sine = 16'h59f3;
    11'd771: sine = 16'h59ab;
    11'd772: sine = 16'h5963;
    11'd773: sine = 16'h591b;
    11'd774: sine = 16'h58d3;
    11'd775: sine = 16'h588a;
    11'd776: sine = 16'h5842;
    11'd777: sine = 16'h57f9;
    11'd778: sine = 16'h57b0;
    11'd779: sine = 16'h5766;
    11'd780: sine = 16'h571d;
    11'd781: sine = 16'h56d3;
    11'd782: sine = 16'h5689;
    11'd783: sine = 16'h563f;
    11'd784: sine = 16'h55f4;
    11'd785: sine = 16'h55aa;
    11'd786: sine = 16'h555f;
    11'd787: sine = 16'h5514;
    11'd788: sine = 16'h54c9;
    11'd789: sine = 16'h547d;
    11'd790: sine = 16'h5432;
    11'd791: sine = 16'h53e6;
    11'd792: sine = 16'h539a;
    11'd793: sine = 16'h534e;
    11'd794: sine = 16'h5301;
    11'd795: sine = 16'h52b5;
    11'd796: sine = 16'h5268;
    11'd797: sine = 16'h521b;
    11'd798: sine = 16'h51ce;
    11'd799: sine = 16'h5180;
    11'd800: sine = 16'h5133;
    11'd801: sine = 16'h50e5;
    11'd802: sine = 16'h5097;
    11'd803: sine = 16'h5049;
    11'd804: sine = 16'h4ffa;
    11'd805: sine = 16'h4fac;
    11'd806: sine = 16'h4f5d;
    11'd807: sine = 16'h4f0e;
    11'd808: sine = 16'h4ebf;
    11'd809: sine = 16'h4e6f;
    11'd810: sine = 16'h4e20;
    11'd811: sine = 16'h4dd0;
    11'd812: sine = 16'h4d80;
    11'd813: sine = 16'h4d30;
    11'd814: sine = 16'h4ce0;
    11'd815: sine = 16'h4c8f;
    11'd816: sine = 16'h4c3f;
    11'd817: sine = 16'h4bee;
    11'd818: sine = 16'h4b9d;
    11'd819: sine = 16'h4b4c;
    11'd820: sine = 16'h4afa;
    11'd821: sine = 16'h4aa9;
    11'd822: sine = 16'h4a57;
    11'd823: sine = 16'h4a05;
    11'd824: sine = 16'h49b3;
    11'd825: sine = 16'h4961;
    11'd826: sine = 16'h490e;
    11'd827: sine = 16'h48bc;
    11'd828: sine = 16'h4869;
    11'd829: sine = 16'h4816;
    11'd830: sine = 16'h47c3;
    11'd831: sine = 16'h476f;
    11'd832: sine = 16'h471c;
    11'd833: sine = 16'h46c8;
    11'd834: sine = 16'h4674;
    11'd835: sine = 16'h4620;
    11'd836: sine = 16'h45cc;
    11'd837: sine = 16'h4578;
    11'd838: sine = 16'h4523;
    11'd839: sine = 16'h44cf;
    11'd840: sine = 16'h447a;
    11'd841: sine = 16'h4425;
    11'd842: sine = 16'h43d0;
    11'd843: sine = 16'h437a;
    11'd844: sine = 16'h4325;
    11'd845: sine = 16'h42cf;
    11'd846: sine = 16'h4279;
    11'd847: sine = 16'h4223;
    11'd848: sine = 16'h41cd;
    11'd849: sine = 16'h4177;
    11'd850: sine = 16'h4120;
    11'd851: sine = 16'h40ca;
    11'd852: sine = 16'h4073;
    11'd853: sine = 16'h401c;
    11'd854: sine = 16'h3fc5;
    11'd855: sine = 16'h3f6e;
    11'd856: sine = 16'h3f16;
    11'd857: sine = 16'h3ebf;
    11'd858: sine = 16'h3e67;
    11'd859: sine = 16'h3e0f;
    11'd860: sine = 16'h3db7;
    11'd861: sine = 16'h3d5f;
    11'd862: sine = 16'h3d07;
    11'd863: sine = 16'h3cae;
    11'd864: sine = 16'h3c56;
    11'd865: sine = 16'h3bfd;
    11'd866: sine = 16'h3ba4;
    11'd867: sine = 16'h3b4b;
    11'd868: sine = 16'h3af2;
    11'd869: sine = 16'h3a99;
    11'd870: sine = 16'h3a3f;
    11'd871: sine = 16'h39e6;
    11'd872: sine = 16'h398c;
    11'd873: sine = 16'h3932;
    11'd874: sine = 16'h38d8;
    11'd875: sine = 16'h387e;
    11'd876: sine = 16'h3824;
    11'd877: sine = 16'h37c9;
    11'd878: sine = 16'h376f;
    11'd879: sine = 16'h3714;
    11'd880: sine = 16'h36b9;
    11'd881: sine = 16'h365e;
    11'd882: sine = 16'h3603;
    11'd883: sine = 16'h35a8;
    11'd884: sine = 16'h354d;
    11'd885: sine = 16'h34f1;
    11'd886: sine = 16'h3496;
    11'd887: sine = 16'h343a;
    11'd888: sine = 16'h33de;
    11'd889: sine = 16'h3382;
    11'd890: sine = 16'h3326;
    11'd891: sine = 16'h32ca;
    11'd892: sine = 16'h326d;
    11'd893: sine = 16'h3211;
    11'd894: sine = 16'h31b4;
    11'd895: sine = 16'h3158;
    11'd896: sine = 16'h30fb;
    11'd897: sine = 16'h309e;
    11'd898: sine = 16'h3041;
    11'd899: sine = 16'h2fe4;
    11'd900: sine = 16'h2f86;
    11'd901: sine = 16'h2f29;
    11'd902: sine = 16'h2ecc;
    11'd903: sine = 16'h2e6e;
    11'd904: sine = 16'h2e10;
    11'd905: sine = 16'h2db2;
    11'd906: sine = 16'h2d54;
    11'd907: sine = 16'h2cf6;
    11'd908: sine = 16'h2c98;
    11'd909: sine = 16'h2c3a;
    11'd910: sine = 16'h2bdb;
    11'd911: sine = 16'h2b7d;
    11'd912: sine = 16'h2b1e;
    11'd913: sine = 16'h2ac0;
    11'd914: sine = 16'h2a61;
    11'd915: sine = 16'h2a02;
    11'd916: sine = 16'h29a3;
    11'd917: sine = 16'h2944;
    11'd918: sine = 16'h28e5;
    11'd919: sine = 16'h2885;
    11'd920: sine = 16'h2826;
    11'd921: sine = 16'h27c6;
    11'd922: sine = 16'h2767;
    11'd923: sine = 16'h2707;
    11'd924: sine = 16'h26a7;
    11'd925: sine = 16'h2647;
    11'd926: sine = 16'h25e7;
    11'd927: sine = 16'h2587;
    11'd928: sine = 16'h2527;
    11'd929: sine = 16'h24c7;
    11'd930: sine = 16'h2467;
    11'd931: sine = 16'h2406;
    11'd932: sine = 16'h23a6;
    11'd933: sine = 16'h2345;
    11'd934: sine = 16'h22e4;
    11'd935: sine = 16'h2284;
    11'd936: sine = 16'h2223;
    11'd937: sine = 16'h21c2;
    11'd938: sine = 16'h2161;
    11'd939: sine = 16'h2100;
    11'd940: sine = 16'h209f;
    11'd941: sine = 16'h203d;
    11'd942: sine = 16'h1fdc;
    11'd943: sine = 16'h1f7b;
    11'd944: sine = 16'h1f19;
    11'd945: sine = 16'h1eb8;
    11'd946: sine = 16'h1e56;
    11'd947: sine = 16'h1df4;
    11'd948: sine = 16'h1d93;
    11'd949: sine = 16'h1d31;
    11'd950: sine = 16'h1ccf;
    11'd951: sine = 16'h1c6d;
    11'd952: sine = 16'h1c0b;
    11'd953: sine = 16'h1ba9;
    11'd954: sine = 16'h1b46;
    11'd955: sine = 16'h1ae4;
    11'd956: sine = 16'h1a82;
    11'd957: sine = 16'h1a20;
    11'd958: sine = 16'h19bd;
    11'd959: sine = 16'h195b;
    11'd960: sine = 16'h18f8;
    11'd961: sine = 16'h1895;
    11'd962: sine = 16'h1833;
    11'd963: sine = 16'h17d0;
    11'd964: sine = 16'h176d;
    11'd965: sine = 16'h170a;
    11'd966: sine = 16'h16a7;
    11'd967: sine = 16'h1644;
    11'd968: sine = 16'h15e1;
    11'd969: sine = 16'h157e;
    11'd970: sine = 16'h151b;
    11'd971: sine = 16'h14b8;
    11'd972: sine = 16'h1455;
    11'd973: sine = 16'h13f2;
    11'd974: sine = 16'h138e;
    11'd975: sine = 16'h132b;
    11'd976: sine = 16'h12c7;
    11'd977: sine = 16'h1264;
    11'd978: sine = 16'h1200;
    11'd979: sine = 16'h119d;
    11'd980: sine = 16'h1139;
    11'd981: sine = 16'h10d6;
    11'd982: sine = 16'h1072;
    11'd983: sine = 16'h100e;
    11'd984: sine = 16'hfab;
    11'd985: sine = 16'hf47;
    11'd986: sine = 16'hee3;
    11'd987: sine = 16'he7f;
    11'd988: sine = 16'he1b;
    11'd989: sine = 16'hdb7;
    11'd990: sine = 16'hd53;
    11'd991: sine = 16'hcef;
    11'd992: sine = 16'hc8b;
    11'd993: sine = 16'hc27;
    11'd994: sine = 16'hbc3;
    11'd995: sine = 16'hb5f;
    11'd996: sine = 16'hafb;
    11'd997: sine = 16'ha97;
    11'd998: sine = 16'ha32;
    11'd999: sine = 16'h9ce;
    11'd1000: sine = 16'h96a;
    11'd1001: sine = 16'h906;
    11'd1002: sine = 16'h8a1;
    11'd1003: sine = 16'h83d;
    11'd1004: sine = 16'h7d9;
    11'd1005: sine = 16'h774;
    11'd1006: sine = 16'h710;
    11'd1007: sine = 16'h6ac;
    11'd1008: sine = 16'h647;
    11'd1009: sine = 16'h5e3;
    11'd1010: sine = 16'h57e;
    11'd1011: sine = 16'h51a;
    11'd1012: sine = 16'h4b6;
    11'd1013: sine = 16'h451;
    11'd1014: sine = 16'h3ed;
    11'd1015: sine = 16'h388;
    11'd1016: sine = 16'h324;
    11'd1017: sine = 16'h2bf;
    11'd1018: sine = 16'h25b;
    11'd1019: sine = 16'h1f6;
    11'd1020: sine = 16'h192;
    11'd1021: sine = 16'h12d;
    11'd1022: sine = 16'hc9;
    11'd1023: sine = 16'h64;
    11'd1024: sine = 16'h0;
    11'd1025: sine = 16'hff9c;
    11'd1026: sine = 16'hff37;
    11'd1027: sine = 16'hfed3;
    11'd1028: sine = 16'hfe6e;
    11'd1029: sine = 16'hfe0a;
    11'd1030: sine = 16'hfda5;
    11'd1031: sine = 16'hfd41;
    11'd1032: sine = 16'hfcdc;
    11'd1033: sine = 16'hfc78;
    11'd1034: sine = 16'hfc13;
    11'd1035: sine = 16'hfbaf;
    11'd1036: sine = 16'hfb4a;
    11'd1037: sine = 16'hfae6;
    11'd1038: sine = 16'hfa82;
    11'd1039: sine = 16'hfa1d;
    11'd1040: sine = 16'hf9b9;
    11'd1041: sine = 16'hf954;
    11'd1042: sine = 16'hf8f0;
    11'd1043: sine = 16'hf88c;
    11'd1044: sine = 16'hf827;
    11'd1045: sine = 16'hf7c3;
    11'd1046: sine = 16'hf75f;
    11'd1047: sine = 16'hf6fa;
    11'd1048: sine = 16'hf696;
    11'd1049: sine = 16'hf632;
    11'd1050: sine = 16'hf5ce;
    11'd1051: sine = 16'hf569;
    11'd1052: sine = 16'hf505;
    11'd1053: sine = 16'hf4a1;
    11'd1054: sine = 16'hf43d;
    11'd1055: sine = 16'hf3d9;
    11'd1056: sine = 16'hf375;
    11'd1057: sine = 16'hf311;
    11'd1058: sine = 16'hf2ad;
    11'd1059: sine = 16'hf249;
    11'd1060: sine = 16'hf1e5;
    11'd1061: sine = 16'hf181;
    11'd1062: sine = 16'hf11d;
    11'd1063: sine = 16'hf0b9;
    11'd1064: sine = 16'hf055;
    11'd1065: sine = 16'heff2;
    11'd1066: sine = 16'hef8e;
    11'd1067: sine = 16'hef2a;
    11'd1068: sine = 16'heec7;
    11'd1069: sine = 16'hee63;
    11'd1070: sine = 16'hee00;
    11'd1071: sine = 16'hed9c;
    11'd1072: sine = 16'hed39;
    11'd1073: sine = 16'hecd5;
    11'd1074: sine = 16'hec72;
    11'd1075: sine = 16'hec0e;
    11'd1076: sine = 16'hebab;
    11'd1077: sine = 16'heb48;
    11'd1078: sine = 16'heae5;
    11'd1079: sine = 16'hea82;
    11'd1080: sine = 16'hea1f;
    11'd1081: sine = 16'he9bc;
    11'd1082: sine = 16'he959;
    11'd1083: sine = 16'he8f6;
    11'd1084: sine = 16'he893;
    11'd1085: sine = 16'he830;
    11'd1086: sine = 16'he7cd;
    11'd1087: sine = 16'he76b;
    11'd1088: sine = 16'he708;
    11'd1089: sine = 16'he6a5;
    11'd1090: sine = 16'he643;
    11'd1091: sine = 16'he5e0;
    11'd1092: sine = 16'he57e;
    11'd1093: sine = 16'he51c;
    11'd1094: sine = 16'he4ba;
    11'd1095: sine = 16'he457;
    11'd1096: sine = 16'he3f5;
    11'd1097: sine = 16'he393;
    11'd1098: sine = 16'he331;
    11'd1099: sine = 16'he2cf;
    11'd1100: sine = 16'he26d;
    11'd1101: sine = 16'he20c;
    11'd1102: sine = 16'he1aa;
    11'd1103: sine = 16'he148;
    11'd1104: sine = 16'he0e7;
    11'd1105: sine = 16'he085;
    11'd1106: sine = 16'he024;
    11'd1107: sine = 16'hdfc3;
    11'd1108: sine = 16'hdf61;
    11'd1109: sine = 16'hdf00;
    11'd1110: sine = 16'hde9f;
    11'd1111: sine = 16'hde3e;
    11'd1112: sine = 16'hdddd;
    11'd1113: sine = 16'hdd7c;
    11'd1114: sine = 16'hdd1c;
    11'd1115: sine = 16'hdcbb;
    11'd1116: sine = 16'hdc5a;
    11'd1117: sine = 16'hdbfa;
    11'd1118: sine = 16'hdb99;
    11'd1119: sine = 16'hdb39;
    11'd1120: sine = 16'hdad9;
    11'd1121: sine = 16'hda79;
    11'd1122: sine = 16'hda19;
    11'd1123: sine = 16'hd9b9;
    11'd1124: sine = 16'hd959;
    11'd1125: sine = 16'hd8f9;
    11'd1126: sine = 16'hd899;
    11'd1127: sine = 16'hd83a;
    11'd1128: sine = 16'hd7da;
    11'd1129: sine = 16'hd77b;
    11'd1130: sine = 16'hd71b;
    11'd1131: sine = 16'hd6bc;
    11'd1132: sine = 16'hd65d;
    11'd1133: sine = 16'hd5fe;
    11'd1134: sine = 16'hd59f;
    11'd1135: sine = 16'hd540;
    11'd1136: sine = 16'hd4e2;
    11'd1137: sine = 16'hd483;
    11'd1138: sine = 16'hd425;
    11'd1139: sine = 16'hd3c6;
    11'd1140: sine = 16'hd368;
    11'd1141: sine = 16'hd30a;
    11'd1142: sine = 16'hd2ac;
    11'd1143: sine = 16'hd24e;
    11'd1144: sine = 16'hd1f0;
    11'd1145: sine = 16'hd192;
    11'd1146: sine = 16'hd134;
    11'd1147: sine = 16'hd0d7;
    11'd1148: sine = 16'hd07a;
    11'd1149: sine = 16'hd01c;
    11'd1150: sine = 16'hcfbf;
    11'd1151: sine = 16'hcf62;
    11'd1152: sine = 16'hcf05;
    11'd1153: sine = 16'hcea8;
    11'd1154: sine = 16'hce4c;
    11'd1155: sine = 16'hcdef;
    11'd1156: sine = 16'hcd93;
    11'd1157: sine = 16'hcd36;
    11'd1158: sine = 16'hccda;
    11'd1159: sine = 16'hcc7e;
    11'd1160: sine = 16'hcc22;
    11'd1161: sine = 16'hcbc6;
    11'd1162: sine = 16'hcb6a;
    11'd1163: sine = 16'hcb0f;
    11'd1164: sine = 16'hcab3;
    11'd1165: sine = 16'hca58;
    11'd1166: sine = 16'hc9fd;
    11'd1167: sine = 16'hc9a2;
    11'd1168: sine = 16'hc947;
    11'd1169: sine = 16'hc8ec;
    11'd1170: sine = 16'hc891;
    11'd1171: sine = 16'hc837;
    11'd1172: sine = 16'hc7dc;
    11'd1173: sine = 16'hc782;
    11'd1174: sine = 16'hc728;
    11'd1175: sine = 16'hc6ce;
    11'd1176: sine = 16'hc674;
    11'd1177: sine = 16'hc61a;
    11'd1178: sine = 16'hc5c1;
    11'd1179: sine = 16'hc567;
    11'd1180: sine = 16'hc50e;
    11'd1181: sine = 16'hc4b5;
    11'd1182: sine = 16'hc45c;
    11'd1183: sine = 16'hc403;
    11'd1184: sine = 16'hc3aa;
    11'd1185: sine = 16'hc352;
    11'd1186: sine = 16'hc2f9;
    11'd1187: sine = 16'hc2a1;
    11'd1188: sine = 16'hc249;
    11'd1189: sine = 16'hc1f1;
    11'd1190: sine = 16'hc199;
    11'd1191: sine = 16'hc141;
    11'd1192: sine = 16'hc0ea;
    11'd1193: sine = 16'hc092;
    11'd1194: sine = 16'hc03b;
    11'd1195: sine = 16'hbfe4;
    11'd1196: sine = 16'hbf8d;
    11'd1197: sine = 16'hbf36;
    11'd1198: sine = 16'hbee0;
    11'd1199: sine = 16'hbe89;
    11'd1200: sine = 16'hbe33;
    11'd1201: sine = 16'hbddd;
    11'd1202: sine = 16'hbd87;
    11'd1203: sine = 16'hbd31;
    11'd1204: sine = 16'hbcdb;
    11'd1205: sine = 16'hbc86;
    11'd1206: sine = 16'hbc30;
    11'd1207: sine = 16'hbbdb;
    11'd1208: sine = 16'hbb86;
    11'd1209: sine = 16'hbb31;
    11'd1210: sine = 16'hbadd;
    11'd1211: sine = 16'hba88;
    11'd1212: sine = 16'hba34;
    11'd1213: sine = 16'hb9e0;
    11'd1214: sine = 16'hb98c;
    11'd1215: sine = 16'hb938;
    11'd1216: sine = 16'hb8e4;
    11'd1217: sine = 16'hb891;
    11'd1218: sine = 16'hb83d;
    11'd1219: sine = 16'hb7ea;
    11'd1220: sine = 16'hb797;
    11'd1221: sine = 16'hb744;
    11'd1222: sine = 16'hb6f2;
    11'd1223: sine = 16'hb69f;
    11'd1224: sine = 16'hb64d;
    11'd1225: sine = 16'hb5fb;
    11'd1226: sine = 16'hb5a9;
    11'd1227: sine = 16'hb557;
    11'd1228: sine = 16'hb506;
    11'd1229: sine = 16'hb4b4;
    11'd1230: sine = 16'hb463;
    11'd1231: sine = 16'hb412;
    11'd1232: sine = 16'hb3c1;
    11'd1233: sine = 16'hb371;
    11'd1234: sine = 16'hb320;
    11'd1235: sine = 16'hb2d0;
    11'd1236: sine = 16'hb280;
    11'd1237: sine = 16'hb230;
    11'd1238: sine = 16'hb1e0;
    11'd1239: sine = 16'hb191;
    11'd1240: sine = 16'hb141;
    11'd1241: sine = 16'hb0f2;
    11'd1242: sine = 16'hb0a3;
    11'd1243: sine = 16'hb054;
    11'd1244: sine = 16'hb006;
    11'd1245: sine = 16'hafb7;
    11'd1246: sine = 16'haf69;
    11'd1247: sine = 16'haf1b;
    11'd1248: sine = 16'haecd;
    11'd1249: sine = 16'hae80;
    11'd1250: sine = 16'hae32;
    11'd1251: sine = 16'hade5;
    11'd1252: sine = 16'had98;
    11'd1253: sine = 16'had4b;
    11'd1254: sine = 16'hacff;
    11'd1255: sine = 16'hacb2;
    11'd1256: sine = 16'hac66;
    11'd1257: sine = 16'hac1a;
    11'd1258: sine = 16'habce;
    11'd1259: sine = 16'hab83;
    11'd1260: sine = 16'hab37;
    11'd1261: sine = 16'haaec;
    11'd1262: sine = 16'haaa1;
    11'd1263: sine = 16'haa56;
    11'd1264: sine = 16'haa0c;
    11'd1265: sine = 16'ha9c1;
    11'd1266: sine = 16'ha977;
    11'd1267: sine = 16'ha92d;
    11'd1268: sine = 16'ha8e3;
    11'd1269: sine = 16'ha89a;
    11'd1270: sine = 16'ha850;
    11'd1271: sine = 16'ha807;
    11'd1272: sine = 16'ha7be;
    11'd1273: sine = 16'ha776;
    11'd1274: sine = 16'ha72d;
    11'd1275: sine = 16'ha6e5;
    11'd1276: sine = 16'ha69d;
    11'd1277: sine = 16'ha655;
    11'd1278: sine = 16'ha60d;
    11'd1279: sine = 16'ha5c6;
    11'd1280: sine = 16'ha57f;
    11'd1281: sine = 16'ha538;
    11'd1282: sine = 16'ha4f1;
    11'd1283: sine = 16'ha4aa;
    11'd1284: sine = 16'ha464;
    11'd1285: sine = 16'ha41e;
    11'd1286: sine = 16'ha3d8;
    11'd1287: sine = 16'ha393;
    11'd1288: sine = 16'ha34d;
    11'd1289: sine = 16'ha308;
    11'd1290: sine = 16'ha2c3;
    11'd1291: sine = 16'ha27e;
    11'd1292: sine = 16'ha23a;
    11'd1293: sine = 16'ha1f5;
    11'd1294: sine = 16'ha1b1;
    11'd1295: sine = 16'ha16d;
    11'd1296: sine = 16'ha12a;
    11'd1297: sine = 16'ha0e6;
    11'd1298: sine = 16'ha0a3;
    11'd1299: sine = 16'ha060;
    11'd1300: sine = 16'ha01e;
    11'd1301: sine = 16'h9fdb;
    11'd1302: sine = 16'h9f99;
    11'd1303: sine = 16'h9f57;
    11'd1304: sine = 16'h9f15;
    11'd1305: sine = 16'h9ed3;
    11'd1306: sine = 16'h9e92;
    11'd1307: sine = 16'h9e51;
    11'd1308: sine = 16'h9e10;
    11'd1309: sine = 16'h9dd0;
    11'd1310: sine = 16'h9d8f;
    11'd1311: sine = 16'h9d4f;
    11'd1312: sine = 16'h9d0f;
    11'd1313: sine = 16'h9cd0;
    11'd1314: sine = 16'h9c90;
    11'd1315: sine = 16'h9c51;
    11'd1316: sine = 16'h9c12;
    11'd1317: sine = 16'h9bd3;
    11'd1318: sine = 16'h9b95;
    11'd1319: sine = 16'h9b57;
    11'd1320: sine = 16'h9b19;
    11'd1321: sine = 16'h9adb;
    11'd1322: sine = 16'h9a9e;
    11'd1323: sine = 16'h9a60;
    11'd1324: sine = 16'h9a23;
    11'd1325: sine = 16'h99e7;
    11'd1326: sine = 16'h99aa;
    11'd1327: sine = 16'h996e;
    11'd1328: sine = 16'h9932;
    11'd1329: sine = 16'h98f6;
    11'd1330: sine = 16'h98bb;
    11'd1331: sine = 16'h987f;
    11'd1332: sine = 16'h9844;
    11'd1333: sine = 16'h9809;
    11'd1334: sine = 16'h97cf;
    11'd1335: sine = 16'h9795;
    11'd1336: sine = 16'h975b;
    11'd1337: sine = 16'h9721;
    11'd1338: sine = 16'h96e7;
    11'd1339: sine = 16'h96ae;
    11'd1340: sine = 16'h9675;
    11'd1341: sine = 16'h963c;
    11'd1342: sine = 16'h9604;
    11'd1343: sine = 16'h95cc;
    11'd1344: sine = 16'h9594;
    11'd1345: sine = 16'h955c;
    11'd1346: sine = 16'h9525;
    11'd1347: sine = 16'h94ed;
    11'd1348: sine = 16'h94b6;
    11'd1349: sine = 16'h9480;
    11'd1350: sine = 16'h9449;
    11'd1351: sine = 16'h9413;
    11'd1352: sine = 16'h93dd;
    11'd1353: sine = 16'h93a8;
    11'd1354: sine = 16'h9372;
    11'd1355: sine = 16'h933d;
    11'd1356: sine = 16'h9308;
    11'd1357: sine = 16'h92d4;
    11'd1358: sine = 16'h929f;
    11'd1359: sine = 16'h926b;
    11'd1360: sine = 16'h9237;
    11'd1361: sine = 16'h9204;
    11'd1362: sine = 16'h91d0;
    11'd1363: sine = 16'h919d;
    11'd1364: sine = 16'h916b;
    11'd1365: sine = 16'h9138;
    11'd1366: sine = 16'h9106;
    11'd1367: sine = 16'h90d4;
    11'd1368: sine = 16'h90a2;
    11'd1369: sine = 16'h9071;
    11'd1370: sine = 16'h9040;
    11'd1371: sine = 16'h900f;
    11'd1372: sine = 16'h8fde;
    11'd1373: sine = 16'h8fae;
    11'd1374: sine = 16'h8f7e;
    11'd1375: sine = 16'h8f4e;
    11'd1376: sine = 16'h8f1f;
    11'd1377: sine = 16'h8eef;
    11'd1378: sine = 16'h8ec0;
    11'd1379: sine = 16'h8e92;
    11'd1380: sine = 16'h8e63;
    11'd1381: sine = 16'h8e35;
    11'd1382: sine = 16'h8e07;
    11'd1383: sine = 16'h8dda;
    11'd1384: sine = 16'h8dac;
    11'd1385: sine = 16'h8d7f;
    11'd1386: sine = 16'h8d52;
    11'd1387: sine = 16'h8d26;
    11'd1388: sine = 16'h8cfa;
    11'd1389: sine = 16'h8cce;
    11'd1390: sine = 16'h8ca2;
    11'd1391: sine = 16'h8c77;
    11'd1392: sine = 16'h8c4b;
    11'd1393: sine = 16'h8c21;
    11'd1394: sine = 16'h8bf6;
    11'd1395: sine = 16'h8bcc;
    11'd1396: sine = 16'h8ba2;
    11'd1397: sine = 16'h8b78;
    11'd1398: sine = 16'h8b4f;
    11'd1399: sine = 16'h8b25;
    11'd1400: sine = 16'h8afd;
    11'd1401: sine = 16'h8ad4;
    11'd1402: sine = 16'h8aac;
    11'd1403: sine = 16'h8a84;
    11'd1404: sine = 16'h8a5c;
    11'd1405: sine = 16'h8a34;
    11'd1406: sine = 16'h8a0d;
    11'd1407: sine = 16'h89e6;
    11'd1408: sine = 16'h89c0;
    11'd1409: sine = 16'h8999;
    11'd1410: sine = 16'h8973;
    11'd1411: sine = 16'h894e;
    11'd1412: sine = 16'h8928;
    11'd1413: sine = 16'h8903;
    11'd1414: sine = 16'h88de;
    11'd1415: sine = 16'h88b9;
    11'd1416: sine = 16'h8895;
    11'd1417: sine = 16'h8871;
    11'd1418: sine = 16'h884d;
    11'd1419: sine = 16'h882a;
    11'd1420: sine = 16'h8807;
    11'd1421: sine = 16'h87e4;
    11'd1422: sine = 16'h87c1;
    11'd1423: sine = 16'h879f;
    11'd1424: sine = 16'h877d;
    11'd1425: sine = 16'h875b;
    11'd1426: sine = 16'h873a;
    11'd1427: sine = 16'h8719;
    11'd1428: sine = 16'h86f8;
    11'd1429: sine = 16'h86d7;
    11'd1430: sine = 16'h86b7;
    11'd1431: sine = 16'h8697;
    11'd1432: sine = 16'h8677;
    11'd1433: sine = 16'h8658;
    11'd1434: sine = 16'h8639;
    11'd1435: sine = 16'h861a;
    11'd1436: sine = 16'h85fc;
    11'd1437: sine = 16'h85dd;
    11'd1438: sine = 16'h85bf;
    11'd1439: sine = 16'h85a2;
    11'd1440: sine = 16'h8584;
    11'd1441: sine = 16'h8567;
    11'd1442: sine = 16'h854b;
    11'd1443: sine = 16'h852e;
    11'd1444: sine = 16'h8512;
    11'd1445: sine = 16'h84f6;
    11'd1446: sine = 16'h84db;
    11'd1447: sine = 16'h84bf;
    11'd1448: sine = 16'h84a4;
    11'd1449: sine = 16'h848a;
    11'd1450: sine = 16'h846f;
    11'd1451: sine = 16'h8455;
    11'd1452: sine = 16'h843c;
    11'd1453: sine = 16'h8422;
    11'd1454: sine = 16'h8409;
    11'd1455: sine = 16'h83f0;
    11'd1456: sine = 16'h83d7;
    11'd1457: sine = 16'h83bf;
    11'd1458: sine = 16'h83a7;
    11'd1459: sine = 16'h8390;
    11'd1460: sine = 16'h8378;
    11'd1461: sine = 16'h8361;
    11'd1462: sine = 16'h834a;
    11'd1463: sine = 16'h8334;
    11'd1464: sine = 16'h831e;
    11'd1465: sine = 16'h8308;
    11'd1466: sine = 16'h82f2;
    11'd1467: sine = 16'h82dd;
    11'd1468: sine = 16'h82c8;
    11'd1469: sine = 16'h82b3;
    11'd1470: sine = 16'h829f;
    11'd1471: sine = 16'h828b;
    11'd1472: sine = 16'h8277;
    11'd1473: sine = 16'h8264;
    11'd1474: sine = 16'h8250;
    11'd1475: sine = 16'h823e;
    11'd1476: sine = 16'h822b;
    11'd1477: sine = 16'h8219;
    11'd1478: sine = 16'h8207;
    11'd1479: sine = 16'h81f5;
    11'd1480: sine = 16'h81e4;
    11'd1481: sine = 16'h81d3;
    11'd1482: sine = 16'h81c2;
    11'd1483: sine = 16'h81b2;
    11'd1484: sine = 16'h81a2;
    11'd1485: sine = 16'h8192;
    11'd1486: sine = 16'h8182;
    11'd1487: sine = 16'h8173;
    11'd1488: sine = 16'h8164;
    11'd1489: sine = 16'h8156;
    11'd1490: sine = 16'h8147;
    11'd1491: sine = 16'h8139;
    11'd1492: sine = 16'h812c;
    11'd1493: sine = 16'h811e;
    11'd1494: sine = 16'h8111;
    11'd1495: sine = 16'h8104;
    11'd1496: sine = 16'h80f8;
    11'd1497: sine = 16'h80ec;
    11'd1498: sine = 16'h80e0;
    11'd1499: sine = 16'h80d4;
    11'd1500: sine = 16'h80c9;
    11'd1501: sine = 16'h80be;
    11'd1502: sine = 16'h80b4;
    11'd1503: sine = 16'h80a9;
    11'd1504: sine = 16'h809f;
    11'd1505: sine = 16'h8096;
    11'd1506: sine = 16'h808c;
    11'd1507: sine = 16'h8083;
    11'd1508: sine = 16'h807a;
    11'd1509: sine = 16'h8072;
    11'd1510: sine = 16'h806a;
    11'd1511: sine = 16'h8062;
    11'd1512: sine = 16'h805a;
    11'd1513: sine = 16'h8053;
    11'd1514: sine = 16'h804c;
    11'd1515: sine = 16'h8045;
    11'd1516: sine = 16'h803f;
    11'd1517: sine = 16'h8039;
    11'd1518: sine = 16'h8033;
    11'd1519: sine = 16'h802e;
    11'd1520: sine = 16'h8029;
    11'd1521: sine = 16'h8024;
    11'd1522: sine = 16'h8020;
    11'd1523: sine = 16'h801c;
    11'd1524: sine = 16'h8018;
    11'd1525: sine = 16'h8014;
    11'd1526: sine = 16'h8011;
    11'd1527: sine = 16'h800e;
    11'd1528: sine = 16'h800b;
    11'd1529: sine = 16'h8009;
    11'd1530: sine = 16'h8007;
    11'd1531: sine = 16'h8005;
    11'd1532: sine = 16'h8004;
    11'd1533: sine = 16'h8003;
    11'd1534: sine = 16'h8002;
    11'd1535: sine = 16'h8002;
    11'd1536: sine = 16'h8002;
    11'd1537: sine = 16'h8002;
    11'd1538: sine = 16'h8002;
    11'd1539: sine = 16'h8003;
    11'd1540: sine = 16'h8004;
    11'd1541: sine = 16'h8005;
    11'd1542: sine = 16'h8007;
    11'd1543: sine = 16'h8009;
    11'd1544: sine = 16'h800b;
    11'd1545: sine = 16'h800e;
    11'd1546: sine = 16'h8011;
    11'd1547: sine = 16'h8014;
    11'd1548: sine = 16'h8018;
    11'd1549: sine = 16'h801c;
    11'd1550: sine = 16'h8020;
    11'd1551: sine = 16'h8024;
    11'd1552: sine = 16'h8029;
    11'd1553: sine = 16'h802e;
    11'd1554: sine = 16'h8033;
    11'd1555: sine = 16'h8039;
    11'd1556: sine = 16'h803f;
    11'd1557: sine = 16'h8045;
    11'd1558: sine = 16'h804c;
    11'd1559: sine = 16'h8053;
    11'd1560: sine = 16'h805a;
    11'd1561: sine = 16'h8062;
    11'd1562: sine = 16'h806a;
    11'd1563: sine = 16'h8072;
    11'd1564: sine = 16'h807a;
    11'd1565: sine = 16'h8083;
    11'd1566: sine = 16'h808c;
    11'd1567: sine = 16'h8096;
    11'd1568: sine = 16'h809f;
    11'd1569: sine = 16'h80a9;
    11'd1570: sine = 16'h80b4;
    11'd1571: sine = 16'h80be;
    11'd1572: sine = 16'h80c9;
    11'd1573: sine = 16'h80d4;
    11'd1574: sine = 16'h80e0;
    11'd1575: sine = 16'h80ec;
    11'd1576: sine = 16'h80f8;
    11'd1577: sine = 16'h8104;
    11'd1578: sine = 16'h8111;
    11'd1579: sine = 16'h811e;
    11'd1580: sine = 16'h812c;
    11'd1581: sine = 16'h8139;
    11'd1582: sine = 16'h8147;
    11'd1583: sine = 16'h8156;
    11'd1584: sine = 16'h8164;
    11'd1585: sine = 16'h8173;
    11'd1586: sine = 16'h8182;
    11'd1587: sine = 16'h8192;
    11'd1588: sine = 16'h81a2;
    11'd1589: sine = 16'h81b2;
    11'd1590: sine = 16'h81c2;
    11'd1591: sine = 16'h81d3;
    11'd1592: sine = 16'h81e4;
    11'd1593: sine = 16'h81f5;
    11'd1594: sine = 16'h8207;
    11'd1595: sine = 16'h8219;
    11'd1596: sine = 16'h822b;
    11'd1597: sine = 16'h823e;
    11'd1598: sine = 16'h8250;
    11'd1599: sine = 16'h8264;
    11'd1600: sine = 16'h8277;
    11'd1601: sine = 16'h828b;
    11'd1602: sine = 16'h829f;
    11'd1603: sine = 16'h82b3;
    11'd1604: sine = 16'h82c8;
    11'd1605: sine = 16'h82dd;
    11'd1606: sine = 16'h82f2;
    11'd1607: sine = 16'h8308;
    11'd1608: sine = 16'h831e;
    11'd1609: sine = 16'h8334;
    11'd1610: sine = 16'h834a;
    11'd1611: sine = 16'h8361;
    11'd1612: sine = 16'h8378;
    11'd1613: sine = 16'h8390;
    11'd1614: sine = 16'h83a7;
    11'd1615: sine = 16'h83bf;
    11'd1616: sine = 16'h83d7;
    11'd1617: sine = 16'h83f0;
    11'd1618: sine = 16'h8409;
    11'd1619: sine = 16'h8422;
    11'd1620: sine = 16'h843c;
    11'd1621: sine = 16'h8455;
    11'd1622: sine = 16'h846f;
    11'd1623: sine = 16'h848a;
    11'd1624: sine = 16'h84a4;
    11'd1625: sine = 16'h84bf;
    11'd1626: sine = 16'h84db;
    11'd1627: sine = 16'h84f6;
    11'd1628: sine = 16'h8512;
    11'd1629: sine = 16'h852e;
    11'd1630: sine = 16'h854b;
    11'd1631: sine = 16'h8567;
    11'd1632: sine = 16'h8584;
    11'd1633: sine = 16'h85a2;
    11'd1634: sine = 16'h85bf;
    11'd1635: sine = 16'h85dd;
    11'd1636: sine = 16'h85fc;
    11'd1637: sine = 16'h861a;
    11'd1638: sine = 16'h8639;
    11'd1639: sine = 16'h8658;
    11'd1640: sine = 16'h8677;
    11'd1641: sine = 16'h8697;
    11'd1642: sine = 16'h86b7;
    11'd1643: sine = 16'h86d7;
    11'd1644: sine = 16'h86f8;
    11'd1645: sine = 16'h8719;
    11'd1646: sine = 16'h873a;
    11'd1647: sine = 16'h875b;
    11'd1648: sine = 16'h877d;
    11'd1649: sine = 16'h879f;
    11'd1650: sine = 16'h87c1;
    11'd1651: sine = 16'h87e4;
    11'd1652: sine = 16'h8807;
    11'd1653: sine = 16'h882a;
    11'd1654: sine = 16'h884d;
    11'd1655: sine = 16'h8871;
    11'd1656: sine = 16'h8895;
    11'd1657: sine = 16'h88b9;
    11'd1658: sine = 16'h88de;
    11'd1659: sine = 16'h8903;
    11'd1660: sine = 16'h8928;
    11'd1661: sine = 16'h894e;
    11'd1662: sine = 16'h8973;
    11'd1663: sine = 16'h8999;
    11'd1664: sine = 16'h89c0;
    11'd1665: sine = 16'h89e6;
    11'd1666: sine = 16'h8a0d;
    11'd1667: sine = 16'h8a34;
    11'd1668: sine = 16'h8a5c;
    11'd1669: sine = 16'h8a84;
    11'd1670: sine = 16'h8aac;
    11'd1671: sine = 16'h8ad4;
    11'd1672: sine = 16'h8afd;
    11'd1673: sine = 16'h8b25;
    11'd1674: sine = 16'h8b4f;
    11'd1675: sine = 16'h8b78;
    11'd1676: sine = 16'h8ba2;
    11'd1677: sine = 16'h8bcc;
    11'd1678: sine = 16'h8bf6;
    11'd1679: sine = 16'h8c21;
    11'd1680: sine = 16'h8c4b;
    11'd1681: sine = 16'h8c77;
    11'd1682: sine = 16'h8ca2;
    11'd1683: sine = 16'h8cce;
    11'd1684: sine = 16'h8cfa;
    11'd1685: sine = 16'h8d26;
    11'd1686: sine = 16'h8d52;
    11'd1687: sine = 16'h8d7f;
    11'd1688: sine = 16'h8dac;
    11'd1689: sine = 16'h8dda;
    11'd1690: sine = 16'h8e07;
    11'd1691: sine = 16'h8e35;
    11'd1692: sine = 16'h8e63;
    11'd1693: sine = 16'h8e92;
    11'd1694: sine = 16'h8ec0;
    11'd1695: sine = 16'h8eef;
    11'd1696: sine = 16'h8f1f;
    11'd1697: sine = 16'h8f4e;
    11'd1698: sine = 16'h8f7e;
    11'd1699: sine = 16'h8fae;
    11'd1700: sine = 16'h8fde;
    11'd1701: sine = 16'h900f;
    11'd1702: sine = 16'h9040;
    11'd1703: sine = 16'h9071;
    11'd1704: sine = 16'h90a2;
    11'd1705: sine = 16'h90d4;
    11'd1706: sine = 16'h9106;
    11'd1707: sine = 16'h9138;
    11'd1708: sine = 16'h916b;
    11'd1709: sine = 16'h919d;
    11'd1710: sine = 16'h91d0;
    11'd1711: sine = 16'h9204;
    11'd1712: sine = 16'h9237;
    11'd1713: sine = 16'h926b;
    11'd1714: sine = 16'h929f;
    11'd1715: sine = 16'h92d4;
    11'd1716: sine = 16'h9308;
    11'd1717: sine = 16'h933d;
    11'd1718: sine = 16'h9372;
    11'd1719: sine = 16'h93a8;
    11'd1720: sine = 16'h93dd;
    11'd1721: sine = 16'h9413;
    11'd1722: sine = 16'h9449;
    11'd1723: sine = 16'h9480;
    11'd1724: sine = 16'h94b6;
    11'd1725: sine = 16'h94ed;
    11'd1726: sine = 16'h9525;
    11'd1727: sine = 16'h955c;
    11'd1728: sine = 16'h9594;
    11'd1729: sine = 16'h95cc;
    11'd1730: sine = 16'h9604;
    11'd1731: sine = 16'h963c;
    11'd1732: sine = 16'h9675;
    11'd1733: sine = 16'h96ae;
    11'd1734: sine = 16'h96e7;
    11'd1735: sine = 16'h9721;
    11'd1736: sine = 16'h975b;
    11'd1737: sine = 16'h9795;
    11'd1738: sine = 16'h97cf;
    11'd1739: sine = 16'h9809;
    11'd1740: sine = 16'h9844;
    11'd1741: sine = 16'h987f;
    11'd1742: sine = 16'h98bb;
    11'd1743: sine = 16'h98f6;
    11'd1744: sine = 16'h9932;
    11'd1745: sine = 16'h996e;
    11'd1746: sine = 16'h99aa;
    11'd1747: sine = 16'h99e7;
    11'd1748: sine = 16'h9a23;
    11'd1749: sine = 16'h9a60;
    11'd1750: sine = 16'h9a9e;
    11'd1751: sine = 16'h9adb;
    11'd1752: sine = 16'h9b19;
    11'd1753: sine = 16'h9b57;
    11'd1754: sine = 16'h9b95;
    11'd1755: sine = 16'h9bd3;
    11'd1756: sine = 16'h9c12;
    11'd1757: sine = 16'h9c51;
    11'd1758: sine = 16'h9c90;
    11'd1759: sine = 16'h9cd0;
    11'd1760: sine = 16'h9d0f;
    11'd1761: sine = 16'h9d4f;
    11'd1762: sine = 16'h9d8f;
    11'd1763: sine = 16'h9dd0;
    11'd1764: sine = 16'h9e10;
    11'd1765: sine = 16'h9e51;
    11'd1766: sine = 16'h9e92;
    11'd1767: sine = 16'h9ed3;
    11'd1768: sine = 16'h9f15;
    11'd1769: sine = 16'h9f57;
    11'd1770: sine = 16'h9f99;
    11'd1771: sine = 16'h9fdb;
    11'd1772: sine = 16'ha01e;
    11'd1773: sine = 16'ha060;
    11'd1774: sine = 16'ha0a3;
    11'd1775: sine = 16'ha0e6;
    11'd1776: sine = 16'ha12a;
    11'd1777: sine = 16'ha16d;
    11'd1778: sine = 16'ha1b1;
    11'd1779: sine = 16'ha1f5;
    11'd1780: sine = 16'ha23a;
    11'd1781: sine = 16'ha27e;
    11'd1782: sine = 16'ha2c3;
    11'd1783: sine = 16'ha308;
    11'd1784: sine = 16'ha34d;
    11'd1785: sine = 16'ha393;
    11'd1786: sine = 16'ha3d8;
    11'd1787: sine = 16'ha41e;
    11'd1788: sine = 16'ha464;
    11'd1789: sine = 16'ha4aa;
    11'd1790: sine = 16'ha4f1;
    11'd1791: sine = 16'ha538;
    11'd1792: sine = 16'ha57f;
    11'd1793: sine = 16'ha5c6;
    11'd1794: sine = 16'ha60d;
    11'd1795: sine = 16'ha655;
    11'd1796: sine = 16'ha69d;
    11'd1797: sine = 16'ha6e5;
    11'd1798: sine = 16'ha72d;
    11'd1799: sine = 16'ha776;
    11'd1800: sine = 16'ha7be;
    11'd1801: sine = 16'ha807;
    11'd1802: sine = 16'ha850;
    11'd1803: sine = 16'ha89a;
    11'd1804: sine = 16'ha8e3;
    11'd1805: sine = 16'ha92d;
    11'd1806: sine = 16'ha977;
    11'd1807: sine = 16'ha9c1;
    11'd1808: sine = 16'haa0c;
    11'd1809: sine = 16'haa56;
    11'd1810: sine = 16'haaa1;
    11'd1811: sine = 16'haaec;
    11'd1812: sine = 16'hab37;
    11'd1813: sine = 16'hab83;
    11'd1814: sine = 16'habce;
    11'd1815: sine = 16'hac1a;
    11'd1816: sine = 16'hac66;
    11'd1817: sine = 16'hacb2;
    11'd1818: sine = 16'hacff;
    11'd1819: sine = 16'had4b;
    11'd1820: sine = 16'had98;
    11'd1821: sine = 16'hade5;
    11'd1822: sine = 16'hae32;
    11'd1823: sine = 16'hae80;
    11'd1824: sine = 16'haecd;
    11'd1825: sine = 16'haf1b;
    11'd1826: sine = 16'haf69;
    11'd1827: sine = 16'hafb7;
    11'd1828: sine = 16'hb006;
    11'd1829: sine = 16'hb054;
    11'd1830: sine = 16'hb0a3;
    11'd1831: sine = 16'hb0f2;
    11'd1832: sine = 16'hb141;
    11'd1833: sine = 16'hb191;
    11'd1834: sine = 16'hb1e0;
    11'd1835: sine = 16'hb230;
    11'd1836: sine = 16'hb280;
    11'd1837: sine = 16'hb2d0;
    11'd1838: sine = 16'hb320;
    11'd1839: sine = 16'hb371;
    11'd1840: sine = 16'hb3c1;
    11'd1841: sine = 16'hb412;
    11'd1842: sine = 16'hb463;
    11'd1843: sine = 16'hb4b4;
    11'd1844: sine = 16'hb506;
    11'd1845: sine = 16'hb557;
    11'd1846: sine = 16'hb5a9;
    11'd1847: sine = 16'hb5fb;
    11'd1848: sine = 16'hb64d;
    11'd1849: sine = 16'hb69f;
    11'd1850: sine = 16'hb6f2;
    11'd1851: sine = 16'hb744;
    11'd1852: sine = 16'hb797;
    11'd1853: sine = 16'hb7ea;
    11'd1854: sine = 16'hb83d;
    11'd1855: sine = 16'hb891;
    11'd1856: sine = 16'hb8e4;
    11'd1857: sine = 16'hb938;
    11'd1858: sine = 16'hb98c;
    11'd1859: sine = 16'hb9e0;
    11'd1860: sine = 16'hba34;
    11'd1861: sine = 16'hba88;
    11'd1862: sine = 16'hbadd;
    11'd1863: sine = 16'hbb31;
    11'd1864: sine = 16'hbb86;
    11'd1865: sine = 16'hbbdb;
    11'd1866: sine = 16'hbc30;
    11'd1867: sine = 16'hbc86;
    11'd1868: sine = 16'hbcdb;
    11'd1869: sine = 16'hbd31;
    11'd1870: sine = 16'hbd87;
    11'd1871: sine = 16'hbddd;
    11'd1872: sine = 16'hbe33;
    11'd1873: sine = 16'hbe89;
    11'd1874: sine = 16'hbee0;
    11'd1875: sine = 16'hbf36;
    11'd1876: sine = 16'hbf8d;
    11'd1877: sine = 16'hbfe4;
    11'd1878: sine = 16'hc03b;
    11'd1879: sine = 16'hc092;
    11'd1880: sine = 16'hc0ea;
    11'd1881: sine = 16'hc141;
    11'd1882: sine = 16'hc199;
    11'd1883: sine = 16'hc1f1;
    11'd1884: sine = 16'hc249;
    11'd1885: sine = 16'hc2a1;
    11'd1886: sine = 16'hc2f9;
    11'd1887: sine = 16'hc352;
    11'd1888: sine = 16'hc3aa;
    11'd1889: sine = 16'hc403;
    11'd1890: sine = 16'hc45c;
    11'd1891: sine = 16'hc4b5;
    11'd1892: sine = 16'hc50e;
    11'd1893: sine = 16'hc567;
    11'd1894: sine = 16'hc5c1;
    11'd1895: sine = 16'hc61a;
    11'd1896: sine = 16'hc674;
    11'd1897: sine = 16'hc6ce;
    11'd1898: sine = 16'hc728;
    11'd1899: sine = 16'hc782;
    11'd1900: sine = 16'hc7dc;
    11'd1901: sine = 16'hc837;
    11'd1902: sine = 16'hc891;
    11'd1903: sine = 16'hc8ec;
    11'd1904: sine = 16'hc947;
    11'd1905: sine = 16'hc9a2;
    11'd1906: sine = 16'hc9fd;
    11'd1907: sine = 16'hca58;
    11'd1908: sine = 16'hcab3;
    11'd1909: sine = 16'hcb0f;
    11'd1910: sine = 16'hcb6a;
    11'd1911: sine = 16'hcbc6;
    11'd1912: sine = 16'hcc22;
    11'd1913: sine = 16'hcc7e;
    11'd1914: sine = 16'hccda;
    11'd1915: sine = 16'hcd36;
    11'd1916: sine = 16'hcd93;
    11'd1917: sine = 16'hcdef;
    11'd1918: sine = 16'hce4c;
    11'd1919: sine = 16'hcea8;
    11'd1920: sine = 16'hcf05;
    11'd1921: sine = 16'hcf62;
    11'd1922: sine = 16'hcfbf;
    11'd1923: sine = 16'hd01c;
    11'd1924: sine = 16'hd07a;
    11'd1925: sine = 16'hd0d7;
    11'd1926: sine = 16'hd134;
    11'd1927: sine = 16'hd192;
    11'd1928: sine = 16'hd1f0;
    11'd1929: sine = 16'hd24e;
    11'd1930: sine = 16'hd2ac;
    11'd1931: sine = 16'hd30a;
    11'd1932: sine = 16'hd368;
    11'd1933: sine = 16'hd3c6;
    11'd1934: sine = 16'hd425;
    11'd1935: sine = 16'hd483;
    11'd1936: sine = 16'hd4e2;
    11'd1937: sine = 16'hd540;
    11'd1938: sine = 16'hd59f;
    11'd1939: sine = 16'hd5fe;
    11'd1940: sine = 16'hd65d;
    11'd1941: sine = 16'hd6bc;
    11'd1942: sine = 16'hd71b;
    11'd1943: sine = 16'hd77b;
    11'd1944: sine = 16'hd7da;
    11'd1945: sine = 16'hd83a;
    11'd1946: sine = 16'hd899;
    11'd1947: sine = 16'hd8f9;
    11'd1948: sine = 16'hd959;
    11'd1949: sine = 16'hd9b9;
    11'd1950: sine = 16'hda19;
    11'd1951: sine = 16'hda79;
    11'd1952: sine = 16'hdad9;
    11'd1953: sine = 16'hdb39;
    11'd1954: sine = 16'hdb99;
    11'd1955: sine = 16'hdbfa;
    11'd1956: sine = 16'hdc5a;
    11'd1957: sine = 16'hdcbb;
    11'd1958: sine = 16'hdd1c;
    11'd1959: sine = 16'hdd7c;
    11'd1960: sine = 16'hdddd;
    11'd1961: sine = 16'hde3e;
    11'd1962: sine = 16'hde9f;
    11'd1963: sine = 16'hdf00;
    11'd1964: sine = 16'hdf61;
    11'd1965: sine = 16'hdfc3;
    11'd1966: sine = 16'he024;
    11'd1967: sine = 16'he085;
    11'd1968: sine = 16'he0e7;
    11'd1969: sine = 16'he148;
    11'd1970: sine = 16'he1aa;
    11'd1971: sine = 16'he20c;
    11'd1972: sine = 16'he26d;
    11'd1973: sine = 16'he2cf;
    11'd1974: sine = 16'he331;
    11'd1975: sine = 16'he393;
    11'd1976: sine = 16'he3f5;
    11'd1977: sine = 16'he457;
    11'd1978: sine = 16'he4ba;
    11'd1979: sine = 16'he51c;
    11'd1980: sine = 16'he57e;
    11'd1981: sine = 16'he5e0;
    11'd1982: sine = 16'he643;
    11'd1983: sine = 16'he6a5;
    11'd1984: sine = 16'he708;
    11'd1985: sine = 16'he76b;
    11'd1986: sine = 16'he7cd;
    11'd1987: sine = 16'he830;
    11'd1988: sine = 16'he893;
    11'd1989: sine = 16'he8f6;
    11'd1990: sine = 16'he959;
    11'd1991: sine = 16'he9bc;
    11'd1992: sine = 16'hea1f;
    11'd1993: sine = 16'hea82;
    11'd1994: sine = 16'heae5;
    11'd1995: sine = 16'heb48;
    11'd1996: sine = 16'hebab;
    11'd1997: sine = 16'hec0e;
    11'd1998: sine = 16'hec72;
    11'd1999: sine = 16'hecd5;
    11'd2000: sine = 16'hed39;
    11'd2001: sine = 16'hed9c;
    11'd2002: sine = 16'hee00;
    11'd2003: sine = 16'hee63;
    11'd2004: sine = 16'heec7;
    11'd2005: sine = 16'hef2a;
    11'd2006: sine = 16'hef8e;
    11'd2007: sine = 16'heff2;
    11'd2008: sine = 16'hf055;
    11'd2009: sine = 16'hf0b9;
    11'd2010: sine = 16'hf11d;
    11'd2011: sine = 16'hf181;
    11'd2012: sine = 16'hf1e5;
    11'd2013: sine = 16'hf249;
    11'd2014: sine = 16'hf2ad;
    11'd2015: sine = 16'hf311;
    11'd2016: sine = 16'hf375;
    11'd2017: sine = 16'hf3d9;
    11'd2018: sine = 16'hf43d;
    11'd2019: sine = 16'hf4a1;
    11'd2020: sine = 16'hf505;
    11'd2021: sine = 16'hf569;
    11'd2022: sine = 16'hf5ce;
    11'd2023: sine = 16'hf632;
    11'd2024: sine = 16'hf696;
    11'd2025: sine = 16'hf6fa;
    11'd2026: sine = 16'hf75f;
    11'd2027: sine = 16'hf7c3;
    11'd2028: sine = 16'hf827;
    11'd2029: sine = 16'hf88c;
    11'd2030: sine = 16'hf8f0;
    11'd2031: sine = 16'hf954;
    11'd2032: sine = 16'hf9b9;
    11'd2033: sine = 16'hfa1d;
    11'd2034: sine = 16'hfa82;
    11'd2035: sine = 16'hfae6;
    11'd2036: sine = 16'hfb4a;
    11'd2037: sine = 16'hfbaf;
    11'd2038: sine = 16'hfc13;
    11'd2039: sine = 16'hfc78;
    11'd2040: sine = 16'hfcdc;
    11'd2041: sine = 16'hfd41;
    11'd2042: sine = 16'hfda5;
    11'd2043: sine = 16'hfe0a;
    11'd2044: sine = 16'hfe6e;
    11'd2045: sine = 16'hfed3;
    11'd2046: sine = 16'hff37;
    11'd2047: sine = 16'hff9c;
  endcase
end
endmodule
