`timescale 1ns/1ns
module sine_table_11bit_float32
(input c,
 input      [10:0] angle,
 output reg [31:0] sine);

always @(posedge c) begin
  case (angle)
    11'd0: sine = 32'h0;
    11'd1: sine = 32'h3b490fc6;
    11'd2: sine = 32'h3bc90f88;
    11'd3: sine = 32'h3c16cb58;
    11'd4: sine = 32'h3c490e90;
    11'd5: sine = 32'h3c7b514b;
    11'd6: sine = 32'h3c96c9b6;
    11'd7: sine = 32'h3cafea69;
    11'd8: sine = 32'h3cc90ab0;
    11'd9: sine = 32'h3ce22a7a;
    11'd10: sine = 32'h3cfb49b9;
    11'd11: sine = 32'h3d0a342f;
    11'd12: sine = 32'h3d16c32c;
    11'd13: sine = 32'h3d2351cb;
    11'd14: sine = 32'h3d2fe006;
    11'd15: sine = 32'h3d3c6dd5;
    11'd16: sine = 32'h3d48fb2f;
    11'd17: sine = 32'h3d55880e;
    11'd18: sine = 32'h3d621468;
    11'd19: sine = 32'h3d6ea038;
    11'd20: sine = 32'h3d7b2b74;
    11'd21: sine = 32'h3d83db0a;
    11'd22: sine = 32'h3d8a2009;
    11'd23: sine = 32'h3d9064b3;
    11'd24: sine = 32'h3d96a904;
    11'd25: sine = 32'h3d9cecf8;
    11'd26: sine = 32'h3da3308c;
    11'd27: sine = 32'h3da973ba;
    11'd28: sine = 32'h3dafb680;
    11'd29: sine = 32'h3db5f8da;
    11'd30: sine = 32'h3dbc3ac3;
    11'd31: sine = 32'h3dc27c38;
    11'd32: sine = 32'h3dc8bd36;
    11'd33: sine = 32'h3dcefdb7;
    11'd34: sine = 32'h3dd53db9;
    11'd35: sine = 32'h3ddb7d37;
    11'd36: sine = 32'h3de1bc2e;
    11'd37: sine = 32'h3de7fa9a;
    11'd38: sine = 32'h3dee3876;
    11'd39: sine = 32'h3df475c0;
    11'd40: sine = 32'h3dfab272;
    11'd41: sine = 32'h3e007745;
    11'd42: sine = 32'h3e039502;
    11'd43: sine = 32'h3e06b26e;
    11'd44: sine = 32'h3e09cf86;
    11'd45: sine = 32'h3e0cec4a;
    11'd46: sine = 32'h3e1008b6;
    11'd47: sine = 32'h3e1324ca;
    11'd48: sine = 32'h3e164083;
    11'd49: sine = 32'h3e195be0;
    11'd50: sine = 32'h3e1c76dd;
    11'd51: sine = 32'h3e1f917b;
    11'd52: sine = 32'h3e22abb5;
    11'd53: sine = 32'h3e25c58c;
    11'd54: sine = 32'h3e28defc;
    11'd55: sine = 32'h3e2bf804;
    11'd56: sine = 32'h3e2f10a2;
    11'd57: sine = 32'h3e3228d4;
    11'd58: sine = 32'h3e354098;
    11'd59: sine = 32'h3e3857ec;
    11'd60: sine = 32'h3e3b6ecf;
    11'd61: sine = 32'h3e3e853e;
    11'd62: sine = 32'h3e419b37;
    11'd63: sine = 32'h3e44b0b9;
    11'd64: sine = 32'h3e47c5c2;
    11'd65: sine = 32'h3e4ada4f;
    11'd66: sine = 32'h3e4dee5f;
    11'd67: sine = 32'h3e5101f1;
    11'd68: sine = 32'h3e541501;
    11'd69: sine = 32'h3e57278e;
    11'd70: sine = 32'h3e5a3997;
    11'd71: sine = 32'h3e5d4b19;
    11'd72: sine = 32'h3e605c13;
    11'd73: sine = 32'h3e636c82;
    11'd74: sine = 32'h3e667c65;
    11'd75: sine = 32'h3e698bba;
    11'd76: sine = 32'h3e6c9a7f;
    11'd77: sine = 32'h3e6fa8b2;
    11'd78: sine = 32'h3e72b651;
    11'd79: sine = 32'h3e75c35a;
    11'd80: sine = 32'h3e78cfcc;
    11'd81: sine = 32'h3e7bdba4;
    11'd82: sine = 32'h3e7ee6e1;
    11'd83: sine = 32'h3e80f8c0;
    11'd84: sine = 32'h3e827dc0;
    11'd85: sine = 32'h3e840270;
    11'd86: sine = 32'h3e8586ce;
    11'd87: sine = 32'h3e870ada;
    11'd88: sine = 32'h3e888e93;
    11'd89: sine = 32'h3e8a11f7;
    11'd90: sine = 32'h3e8b9507;
    11'd91: sine = 32'h3e8d17c0;
    11'd92: sine = 32'h3e8e9a22;
    11'd93: sine = 32'h3e901c2c;
    11'd94: sine = 32'h3e919ddd;
    11'd95: sine = 32'h3e931f35;
    11'd96: sine = 32'h3e94a031;
    11'd97: sine = 32'h3e9620d2;
    11'd98: sine = 32'h3e97a117;
    11'd99: sine = 32'h3e9920fe;
    11'd100: sine = 32'h3e9aa086;
    11'd101: sine = 32'h3e9c1faf;
    11'd102: sine = 32'h3e9d9e78;
    11'd103: sine = 32'h3e9f1cdf;
    11'd104: sine = 32'h3ea09ae4;
    11'd105: sine = 32'h3ea21887;
    11'd106: sine = 32'h3ea395c5;
    11'd107: sine = 32'h3ea5129e;
    11'd108: sine = 32'h3ea68f12;
    11'd109: sine = 32'h3ea80b1f;
    11'd110: sine = 32'h3ea986c4;
    11'd111: sine = 32'h3eab0200;
    11'd112: sine = 32'h3eac7cd3;
    11'd113: sine = 32'h3eadf73c;
    11'd114: sine = 32'h3eaf713a;
    11'd115: sine = 32'h3eb0eacb;
    11'd116: sine = 32'h3eb263ef;
    11'd117: sine = 32'h3eb3dca5;
    11'd118: sine = 32'h3eb554ec;
    11'd119: sine = 32'h3eb6ccc3;
    11'd120: sine = 32'h3eb84429;
    11'd121: sine = 32'h3eb9bb1e;
    11'd122: sine = 32'h3ebb31a0;
    11'd123: sine = 32'h3ebca7af;
    11'd124: sine = 32'h3ebe1d49;
    11'd125: sine = 32'h3ebf926e;
    11'd126: sine = 32'h3ec1071d;
    11'd127: sine = 32'h3ec27b55;
    11'd128: sine = 32'h3ec3ef15;
    11'd129: sine = 32'h3ec5625c;
    11'd130: sine = 32'h3ec6d529;
    11'd131: sine = 32'h3ec8477c;
    11'd132: sine = 32'h3ec9b953;
    11'd133: sine = 32'h3ecb2aae;
    11'd134: sine = 32'h3ecc9b8b;
    11'd135: sine = 32'h3ece0bea;
    11'd136: sine = 32'h3ecf7bca;
    11'd137: sine = 32'h3ed0eb2a;
    11'd138: sine = 32'h3ed25a09;
    11'd139: sine = 32'h3ed3c866;
    11'd140: sine = 32'h3ed53641;
    11'd141: sine = 32'h3ed6a398;
    11'd142: sine = 32'h3ed8106b;
    11'd143: sine = 32'h3ed97cb9;
    11'd144: sine = 32'h3edae880;
    11'd145: sine = 32'h3edc53c0;
    11'd146: sine = 32'h3eddbe79;
    11'd147: sine = 32'h3edf28a9;
    11'd148: sine = 32'h3ee0924f;
    11'd149: sine = 32'h3ee1fb6a;
    11'd150: sine = 32'h3ee363fa;
    11'd151: sine = 32'h3ee4cbfe;
    11'd152: sine = 32'h3ee63375;
    11'd153: sine = 32'h3ee79a5d;
    11'd154: sine = 32'h3ee900b7;
    11'd155: sine = 32'h3eea6681;
    11'd156: sine = 32'h3eebcbbb;
    11'd157: sine = 32'h3eed3063;
    11'd158: sine = 32'h3eee9478;
    11'd159: sine = 32'h3eeff7fb;
    11'd160: sine = 32'h3ef15aea;
    11'd161: sine = 32'h3ef2bd43;
    11'd162: sine = 32'h3ef41f07;
    11'd163: sine = 32'h3ef58034;
    11'd164: sine = 32'h3ef6e0ca;
    11'd165: sine = 32'h3ef840c8;
    11'd166: sine = 32'h3ef9a02c;
    11'd167: sine = 32'h3efafef7;
    11'd168: sine = 32'h3efc5d27;
    11'd169: sine = 32'h3efdbabb;
    11'd170: sine = 32'h3eff17b2;
    11'd171: sine = 32'h3f003a06;
    11'd172: sine = 32'h3f00e7e4;
    11'd173: sine = 32'h3f019573;
    11'd174: sine = 32'h3f0242b1;
    11'd175: sine = 32'h3f02ef9f;
    11'd176: sine = 32'h3f039c3d;
    11'd177: sine = 32'h3f044889;
    11'd178: sine = 32'h3f04f483;
    11'd179: sine = 32'h3f05a02c;
    11'd180: sine = 32'h3f064b82;
    11'd181: sine = 32'h3f06f686;
    11'd182: sine = 32'h3f07a136;
    11'd183: sine = 32'h3f084b92;
    11'd184: sine = 32'h3f08f59a;
    11'd185: sine = 32'h3f099f4e;
    11'd186: sine = 32'h3f0a48ad;
    11'd187: sine = 32'h3f0af1b7;
    11'd188: sine = 32'h3f0b9a6b;
    11'd189: sine = 32'h3f0c42c9;
    11'd190: sine = 32'h3f0cead0;
    11'd191: sine = 32'h3f0d9281;
    11'd192: sine = 32'h3f0e39da;
    11'd193: sine = 32'h3f0ee0db;
    11'd194: sine = 32'h3f0f8784;
    11'd195: sine = 32'h3f102dd5;
    11'd196: sine = 32'h3f10d3cd;
    11'd197: sine = 32'h3f11796b;
    11'd198: sine = 32'h3f121eb0;
    11'd199: sine = 32'h3f12c39a;
    11'd200: sine = 32'h3f13682a;
    11'd201: sine = 32'h3f140c5f;
    11'd202: sine = 32'h3f14b039;
    11'd203: sine = 32'h3f1553b7;
    11'd204: sine = 32'h3f15f6d9;
    11'd205: sine = 32'h3f16999e;
    11'd206: sine = 32'h3f173c07;
    11'd207: sine = 32'h3f17de12;
    11'd208: sine = 32'h3f187fc0;
    11'd209: sine = 32'h3f19210f;
    11'd210: sine = 32'h3f19c200;
    11'd211: sine = 32'h3f1a6292;
    11'd212: sine = 32'h3f1b02c5;
    11'd213: sine = 32'h3f1ba299;
    11'd214: sine = 32'h3f1c420c;
    11'd215: sine = 32'h3f1ce11f;
    11'd216: sine = 32'h3f1d7fd1;
    11'd217: sine = 32'h3f1e1e22;
    11'd218: sine = 32'h3f1ebc12;
    11'd219: sine = 32'h3f1f599f;
    11'd220: sine = 32'h3f1ff6ca;
    11'd221: sine = 32'h3f209393;
    11'd222: sine = 32'h3f212ff9;
    11'd223: sine = 32'h3f21cbfb;
    11'd224: sine = 32'h3f226799;
    11'd225: sine = 32'h3f2302d3;
    11'd226: sine = 32'h3f239da9;
    11'd227: sine = 32'h3f243819;
    11'd228: sine = 32'h3f24d225;
    11'd229: sine = 32'h3f256bca;
    11'd230: sine = 32'h3f26050a;
    11'd231: sine = 32'h3f269de3;
    11'd232: sine = 32'h3f273656;
    11'd233: sine = 32'h3f27ce61;
    11'd234: sine = 32'h3f286605;
    11'd235: sine = 32'h3f28fd41;
    11'd236: sine = 32'h3f299414;
    11'd237: sine = 32'h3f2a2a80;
    11'd238: sine = 32'h3f2ac082;
    11'd239: sine = 32'h3f2b561a;
    11'd240: sine = 32'h3f2beb49;
    11'd241: sine = 32'h3f2c800f;
    11'd242: sine = 32'h3f2d1469;
    11'd243: sine = 32'h3f2da859;
    11'd244: sine = 32'h3f2e3bde;
    11'd245: sine = 32'h3f2ecef7;
    11'd246: sine = 32'h3f2f61a5;
    11'd247: sine = 32'h3f2ff3e6;
    11'd248: sine = 32'h3f3085bb;
    11'd249: sine = 32'h3f311722;
    11'd250: sine = 32'h3f31a81d;
    11'd251: sine = 32'h3f3238aa;
    11'd252: sine = 32'h3f32c8c9;
    11'd253: sine = 32'h3f33587a;
    11'd254: sine = 32'h3f33e7bc;
    11'd255: sine = 32'h3f34768f;
    11'd256: sine = 32'h3f3504f3;
    11'd257: sine = 32'h3f3592e7;
    11'd258: sine = 32'h3f36206b;
    11'd259: sine = 32'h3f36ad7f;
    11'd260: sine = 32'h3f373a22;
    11'd261: sine = 32'h3f37c655;
    11'd262: sine = 32'h3f385215;
    11'd263: sine = 32'h3f38dd65;
    11'd264: sine = 32'h3f396842;
    11'd265: sine = 32'h3f39f2ac;
    11'd266: sine = 32'h3f3a7ca4;
    11'd267: sine = 32'h3f3b0629;
    11'd268: sine = 32'h3f3b8f3b;
    11'd269: sine = 32'h3f3c17d9;
    11'd270: sine = 32'h3f3ca003;
    11'd271: sine = 32'h3f3d27b8;
    11'd272: sine = 32'h3f3daef9;
    11'd273: sine = 32'h3f3e35c5;
    11'd274: sine = 32'h3f3ebc1b;
    11'd275: sine = 32'h3f3f41fc;
    11'd276: sine = 32'h3f3fc767;
    11'd277: sine = 32'h3f404c5c;
    11'd278: sine = 32'h3f40d0d9;
    11'd279: sine = 32'h3f4154e0;
    11'd280: sine = 32'h3f41d870;
    11'd281: sine = 32'h3f425b88;
    11'd282: sine = 32'h3f42de29;
    11'd283: sine = 32'h3f436051;
    11'd284: sine = 32'h3f43e200;
    11'd285: sine = 32'h3f446337;
    11'd286: sine = 32'h3f44e3f5;
    11'd287: sine = 32'h3f456439;
    11'd288: sine = 32'h3f45e403;
    11'd289: sine = 32'h3f466353;
    11'd290: sine = 32'h3f46e229;
    11'd291: sine = 32'h3f476085;
    11'd292: sine = 32'h3f47de65;
    11'd293: sine = 32'h3f485bca;
    11'd294: sine = 32'h3f48d8b3;
    11'd295: sine = 32'h3f495521;
    11'd296: sine = 32'h3f49d112;
    11'd297: sine = 32'h3f4a4c87;
    11'd298: sine = 32'h3f4ac77f;
    11'd299: sine = 32'h3f4b41fa;
    11'd300: sine = 32'h3f4bbbf7;
    11'd301: sine = 32'h3f4c3577;
    11'd302: sine = 32'h3f4cae79;
    11'd303: sine = 32'h3f4d26fd;
    11'd304: sine = 32'h3f4d9f02;
    11'd305: sine = 32'h3f4e1688;
    11'd306: sine = 32'h3f4e8d90;
    11'd307: sine = 32'h3f4f0417;
    11'd308: sine = 32'h3f4f7a1f;
    11'd309: sine = 32'h3f4fefa7;
    11'd310: sine = 32'h3f5064af;
    11'd311: sine = 32'h3f50d936;
    11'd312: sine = 32'h3f514d3d;
    11'd313: sine = 32'h3f51c0c2;
    11'd314: sine = 32'h3f5233c6;
    11'd315: sine = 32'h3f52a648;
    11'd316: sine = 32'h3f531849;
    11'd317: sine = 32'h3f5389c7;
    11'd318: sine = 32'h3f53fac2;
    11'd319: sine = 32'h3f546b3b;
    11'd320: sine = 32'h3f54db31;
    11'd321: sine = 32'h3f554aa4;
    11'd322: sine = 32'h3f55b993;
    11'd323: sine = 32'h3f5627fe;
    11'd324: sine = 32'h3f5695e5;
    11'd325: sine = 32'h3f570347;
    11'd326: sine = 32'h3f577025;
    11'd327: sine = 32'h3f57dc7f;
    11'd328: sine = 32'h3f584853;
    11'd329: sine = 32'h3f58b3a1;
    11'd330: sine = 32'h3f591e6a;
    11'd331: sine = 32'h3f5988ad;
    11'd332: sine = 32'h3f59f26a;
    11'd333: sine = 32'h3f5a5ba0;
    11'd334: sine = 32'h3f5ac450;
    11'd335: sine = 32'h3f5b2c79;
    11'd336: sine = 32'h3f5b941a;
    11'd337: sine = 32'h3f5bfb34;
    11'd338: sine = 32'h3f5c61c6;
    11'd339: sine = 32'h3f5cc7d1;
    11'd340: sine = 32'h3f5d2d53;
    11'd341: sine = 32'h3f5d924d;
    11'd342: sine = 32'h3f5df6be;
    11'd343: sine = 32'h3f5e5aa6;
    11'd344: sine = 32'h3f5ebe05;
    11'd345: sine = 32'h3f5f20db;
    11'd346: sine = 32'h3f5f8327;
    11'd347: sine = 32'h3f5fe4e9;
    11'd348: sine = 32'h3f604621;
    11'd349: sine = 32'h3f60a6cf;
    11'd350: sine = 32'h3f6106f2;
    11'd351: sine = 32'h3f61668a;
    11'd352: sine = 32'h3f61c597;
    11'd353: sine = 32'h3f622419;
    11'd354: sine = 32'h3f628210;
    11'd355: sine = 32'h3f62df7b;
    11'd356: sine = 32'h3f633c59;
    11'd357: sine = 32'h3f6398ac;
    11'd358: sine = 32'h3f63f472;
    11'd359: sine = 32'h3f644fac;
    11'd360: sine = 32'h3f64aa59;
    11'd361: sine = 32'h3f650479;
    11'd362: sine = 32'h3f655e0b;
    11'd363: sine = 32'h3f65b710;
    11'd364: sine = 32'h3f660f87;
    11'd365: sine = 32'h3f666771;
    11'd366: sine = 32'h3f66becc;
    11'd367: sine = 32'h3f671599;
    11'd368: sine = 32'h3f676bd7;
    11'd369: sine = 32'h3f67c187;
    11'd370: sine = 32'h3f6816a8;
    11'd371: sine = 32'h3f686b39;
    11'd372: sine = 32'h3f68bf3b;
    11'd373: sine = 32'h3f6912ae;
    11'd374: sine = 32'h3f696591;
    11'd375: sine = 32'h3f69b7e4;
    11'd376: sine = 32'h3f6a09a6;
    11'd377: sine = 32'h3f6a5ad9;
    11'd378: sine = 32'h3f6aab7a;
    11'd379: sine = 32'h3f6afb8b;
    11'd380: sine = 32'h3f6b4b0b;
    11'd381: sine = 32'h3f6b99fa;
    11'd382: sine = 32'h3f6be858;
    11'd383: sine = 32'h3f6c3624;
    11'd384: sine = 32'h3f6c835e;
    11'd385: sine = 32'h3f6cd007;
    11'd386: sine = 32'h3f6d1c1d;
    11'd387: sine = 32'h3f6d67a1;
    11'd388: sine = 32'h3f6db293;
    11'd389: sine = 32'h3f6dfcf2;
    11'd390: sine = 32'h3f6e46be;
    11'd391: sine = 32'h3f6e8ff7;
    11'd392: sine = 32'h3f6ed89e;
    11'd393: sine = 32'h3f6f20b0;
    11'd394: sine = 32'h3f6f6830;
    11'd395: sine = 32'h3f6faf1b;
    11'd396: sine = 32'h3f6ff573;
    11'd397: sine = 32'h3f703b37;
    11'd398: sine = 32'h3f708066;
    11'd399: sine = 32'h3f70c501;
    11'd400: sine = 32'h3f710908;
    11'd401: sine = 32'h3f714c7a;
    11'd402: sine = 32'h3f718f57;
    11'd403: sine = 32'h3f71d19f;
    11'd404: sine = 32'h3f721352;
    11'd405: sine = 32'h3f725470;
    11'd406: sine = 32'h3f7294f8;
    11'd407: sine = 32'h3f72d4eb;
    11'd408: sine = 32'h3f731447;
    11'd409: sine = 32'h3f73530e;
    11'd410: sine = 32'h3f73913f;
    11'd411: sine = 32'h3f73ced9;
    11'd412: sine = 32'h3f740bdd;
    11'd413: sine = 32'h3f74484b;
    11'd414: sine = 32'h3f748422;
    11'd415: sine = 32'h3f74bf62;
    11'd416: sine = 32'h3f74fa0b;
    11'd417: sine = 32'h3f75341d;
    11'd418: sine = 32'h3f756d97;
    11'd419: sine = 32'h3f75a67a;
    11'd420: sine = 32'h3f75dec6;
    11'd421: sine = 32'h3f76167a;
    11'd422: sine = 32'h3f764d97;
    11'd423: sine = 32'h3f76841b;
    11'd424: sine = 32'h3f76ba07;
    11'd425: sine = 32'h3f76ef5b;
    11'd426: sine = 32'h3f772417;
    11'd427: sine = 32'h3f77583a;
    11'd428: sine = 32'h3f778bc5;
    11'd429: sine = 32'h3f77beb7;
    11'd430: sine = 32'h3f77f110;
    11'd431: sine = 32'h3f7822d1;
    11'd432: sine = 32'h3f7853f8;
    11'd433: sine = 32'h3f788486;
    11'd434: sine = 32'h3f78b47b;
    11'd435: sine = 32'h3f78e3d6;
    11'd436: sine = 32'h3f791298;
    11'd437: sine = 32'h3f7940c0;
    11'd438: sine = 32'h3f796e4e;
    11'd439: sine = 32'h3f799b43;
    11'd440: sine = 32'h3f79c79d;
    11'd441: sine = 32'h3f79f35e;
    11'd442: sine = 32'h3f7a1e84;
    11'd443: sine = 32'h3f7a4910;
    11'd444: sine = 32'h3f7a7302;
    11'd445: sine = 32'h3f7a9c59;
    11'd446: sine = 32'h3f7ac515;
    11'd447: sine = 32'h3f7aed37;
    11'd448: sine = 32'h3f7b14be;
    11'd449: sine = 32'h3f7b3bab;
    11'd450: sine = 32'h3f7b61fc;
    11'd451: sine = 32'h3f7b87b2;
    11'd452: sine = 32'h3f7baccd;
    11'd453: sine = 32'h3f7bd14d;
    11'd454: sine = 32'h3f7bf531;
    11'd455: sine = 32'h3f7c187a;
    11'd456: sine = 32'h3f7c3b28;
    11'd457: sine = 32'h3f7c5d3a;
    11'd458: sine = 32'h3f7c7eb0;
    11'd459: sine = 32'h3f7c9f8a;
    11'd460: sine = 32'h3f7cbfc9;
    11'd461: sine = 32'h3f7cdf6c;
    11'd462: sine = 32'h3f7cfe73;
    11'd463: sine = 32'h3f7d1cdd;
    11'd464: sine = 32'h3f7d3aac;
    11'd465: sine = 32'h3f7d57de;
    11'd466: sine = 32'h3f7d7474;
    11'd467: sine = 32'h3f7d906e;
    11'd468: sine = 32'h3f7dabcb;
    11'd469: sine = 32'h3f7dc68c;
    11'd470: sine = 32'h3f7de0b1;
    11'd471: sine = 32'h3f7dfa38;
    11'd472: sine = 32'h3f7e1323;
    11'd473: sine = 32'h3f7e2b72;
    11'd474: sine = 32'h3f7e4323;
    11'd475: sine = 32'h3f7e5a38;
    11'd476: sine = 32'h3f7e70b0;
    11'd477: sine = 32'h3f7e868b;
    11'd478: sine = 32'h3f7e9bc9;
    11'd479: sine = 32'h3f7eb069;
    11'd480: sine = 32'h3f7ec46d;
    11'd481: sine = 32'h3f7ed7d4;
    11'd482: sine = 32'h3f7eea9d;
    11'd483: sine = 32'h3f7efcc9;
    11'd484: sine = 32'h3f7f0e58;
    11'd485: sine = 32'h3f7f1f49;
    11'd486: sine = 32'h3f7f2f9d;
    11'd487: sine = 32'h3f7f3f54;
    11'd488: sine = 32'h3f7f4e6d;
    11'd489: sine = 32'h3f7f5ce9;
    11'd490: sine = 32'h3f7f6ac7;
    11'd491: sine = 32'h3f7f7808;
    11'd492: sine = 32'h3f7f84ab;
    11'd493: sine = 32'h3f7f90b1;
    11'd494: sine = 32'h3f7f9c18;
    11'd495: sine = 32'h3f7fa6e3;
    11'd496: sine = 32'h3f7fb10f;
    11'd497: sine = 32'h3f7fba9e;
    11'd498: sine = 32'h3f7fc38f;
    11'd499: sine = 32'h3f7fcbe2;
    11'd500: sine = 32'h3f7fd397;
    11'd501: sine = 32'h3f7fdaaf;
    11'd502: sine = 32'h3f7fe129;
    11'd503: sine = 32'h3f7fe705;
    11'd504: sine = 32'h3f7fec43;
    11'd505: sine = 32'h3f7ff0e3;
    11'd506: sine = 32'h3f7ff4e6;
    11'd507: sine = 32'h3f7ff84a;
    11'd508: sine = 32'h3f7ffb11;
    11'd509: sine = 32'h3f7ffd39;
    11'd510: sine = 32'h3f7ffec4;
    11'd511: sine = 32'h3f7fffb1;
    11'd512: sine = 32'h3f800000;
    11'd513: sine = 32'h3f7fffb1;
    11'd514: sine = 32'h3f7ffec4;
    11'd515: sine = 32'h3f7ffd39;
    11'd516: sine = 32'h3f7ffb11;
    11'd517: sine = 32'h3f7ff84a;
    11'd518: sine = 32'h3f7ff4e6;
    11'd519: sine = 32'h3f7ff0e3;
    11'd520: sine = 32'h3f7fec43;
    11'd521: sine = 32'h3f7fe705;
    11'd522: sine = 32'h3f7fe129;
    11'd523: sine = 32'h3f7fdaaf;
    11'd524: sine = 32'h3f7fd398;
    11'd525: sine = 32'h3f7fcbe2;
    11'd526: sine = 32'h3f7fc38f;
    11'd527: sine = 32'h3f7fba9e;
    11'd528: sine = 32'h3f7fb10f;
    11'd529: sine = 32'h3f7fa6e3;
    11'd530: sine = 32'h3f7f9c19;
    11'd531: sine = 32'h3f7f90b1;
    11'd532: sine = 32'h3f7f84ab;
    11'd533: sine = 32'h3f7f7808;
    11'd534: sine = 32'h3f7f6ac7;
    11'd535: sine = 32'h3f7f5ce9;
    11'd536: sine = 32'h3f7f4e6d;
    11'd537: sine = 32'h3f7f3f54;
    11'd538: sine = 32'h3f7f2f9e;
    11'd539: sine = 32'h3f7f1f49;
    11'd540: sine = 32'h3f7f0e58;
    11'd541: sine = 32'h3f7efcc9;
    11'd542: sine = 32'h3f7eea9d;
    11'd543: sine = 32'h3f7ed7d4;
    11'd544: sine = 32'h3f7ec46d;
    11'd545: sine = 32'h3f7eb069;
    11'd546: sine = 32'h3f7e9bc9;
    11'd547: sine = 32'h3f7e868b;
    11'd548: sine = 32'h3f7e70b0;
    11'd549: sine = 32'h3f7e5a38;
    11'd550: sine = 32'h3f7e4323;
    11'd551: sine = 32'h3f7e2b72;
    11'd552: sine = 32'h3f7e1324;
    11'd553: sine = 32'h3f7dfa39;
    11'd554: sine = 32'h3f7de0b1;
    11'd555: sine = 32'h3f7dc68c;
    11'd556: sine = 32'h3f7dabcc;
    11'd557: sine = 32'h3f7d906e;
    11'd558: sine = 32'h3f7d7475;
    11'd559: sine = 32'h3f7d57de;
    11'd560: sine = 32'h3f7d3aac;
    11'd561: sine = 32'h3f7d1cdd;
    11'd562: sine = 32'h3f7cfe73;
    11'd563: sine = 32'h3f7cdf6c;
    11'd564: sine = 32'h3f7cbfc9;
    11'd565: sine = 32'h3f7c9f8b;
    11'd566: sine = 32'h3f7c7eb0;
    11'd567: sine = 32'h3f7c5d3a;
    11'd568: sine = 32'h3f7c3b28;
    11'd569: sine = 32'h3f7c187a;
    11'd570: sine = 32'h3f7bf531;
    11'd571: sine = 32'h3f7bd14d;
    11'd572: sine = 32'h3f7baccd;
    11'd573: sine = 32'h3f7b87b2;
    11'd574: sine = 32'h3f7b61fc;
    11'd575: sine = 32'h3f7b3bab;
    11'd576: sine = 32'h3f7b14bf;
    11'd577: sine = 32'h3f7aed38;
    11'd578: sine = 32'h3f7ac516;
    11'd579: sine = 32'h3f7a9c59;
    11'd580: sine = 32'h3f7a7302;
    11'd581: sine = 32'h3f7a4910;
    11'd582: sine = 32'h3f7a1e84;
    11'd583: sine = 32'h3f79f35e;
    11'd584: sine = 32'h3f79c79d;
    11'd585: sine = 32'h3f799b43;
    11'd586: sine = 32'h3f796e4e;
    11'd587: sine = 32'h3f7940c0;
    11'd588: sine = 32'h3f791298;
    11'd589: sine = 32'h3f78e3d6;
    11'd590: sine = 32'h3f78b47b;
    11'd591: sine = 32'h3f788486;
    11'd592: sine = 32'h3f7853f8;
    11'd593: sine = 32'h3f7822d1;
    11'd594: sine = 32'h3f77f111;
    11'd595: sine = 32'h3f77beb7;
    11'd596: sine = 32'h3f778bc5;
    11'd597: sine = 32'h3f77583b;
    11'd598: sine = 32'h3f772417;
    11'd599: sine = 32'h3f76ef5b;
    11'd600: sine = 32'h3f76ba07;
    11'd601: sine = 32'h3f76841b;
    11'd602: sine = 32'h3f764d97;
    11'd603: sine = 32'h3f76167a;
    11'd604: sine = 32'h3f75dec6;
    11'd605: sine = 32'h3f75a67b;
    11'd606: sine = 32'h3f756d97;
    11'd607: sine = 32'h3f75341d;
    11'd608: sine = 32'h3f74fa0b;
    11'd609: sine = 32'h3f74bf62;
    11'd610: sine = 32'h3f748422;
    11'd611: sine = 32'h3f74484b;
    11'd612: sine = 32'h3f740bde;
    11'd613: sine = 32'h3f73ced9;
    11'd614: sine = 32'h3f73913f;
    11'd615: sine = 32'h3f73530e;
    11'd616: sine = 32'h3f731448;
    11'd617: sine = 32'h3f72d4eb;
    11'd618: sine = 32'h3f7294f8;
    11'd619: sine = 32'h3f725470;
    11'd620: sine = 32'h3f721353;
    11'd621: sine = 32'h3f71d1a0;
    11'd622: sine = 32'h3f718f57;
    11'd623: sine = 32'h3f714c7a;
    11'd624: sine = 32'h3f710908;
    11'd625: sine = 32'h3f70c502;
    11'd626: sine = 32'h3f708067;
    11'd627: sine = 32'h3f703b37;
    11'd628: sine = 32'h3f6ff573;
    11'd629: sine = 32'h3f6faf1c;
    11'd630: sine = 32'h3f6f6830;
    11'd631: sine = 32'h3f6f20b1;
    11'd632: sine = 32'h3f6ed89e;
    11'd633: sine = 32'h3f6e8ff8;
    11'd634: sine = 32'h3f6e46bf;
    11'd635: sine = 32'h3f6dfcf2;
    11'd636: sine = 32'h3f6db293;
    11'd637: sine = 32'h3f6d67a2;
    11'd638: sine = 32'h3f6d1c1e;
    11'd639: sine = 32'h3f6cd007;
    11'd640: sine = 32'h3f6c835f;
    11'd641: sine = 32'h3f6c3624;
    11'd642: sine = 32'h3f6be858;
    11'd643: sine = 32'h3f6b99fb;
    11'd644: sine = 32'h3f6b4b0c;
    11'd645: sine = 32'h3f6afb8c;
    11'd646: sine = 32'h3f6aab7b;
    11'd647: sine = 32'h3f6a5ad9;
    11'd648: sine = 32'h3f6a09a7;
    11'd649: sine = 32'h3f69b7e4;
    11'd650: sine = 32'h3f696591;
    11'd651: sine = 32'h3f6912ae;
    11'd652: sine = 32'h3f68bf3c;
    11'd653: sine = 32'h3f686b3a;
    11'd654: sine = 32'h3f6816a8;
    11'd655: sine = 32'h3f67c188;
    11'd656: sine = 32'h3f676bd8;
    11'd657: sine = 32'h3f671599;
    11'd658: sine = 32'h3f66becd;
    11'd659: sine = 32'h3f666771;
    11'd660: sine = 32'h3f660f88;
    11'd661: sine = 32'h3f65b711;
    11'd662: sine = 32'h3f655e0c;
    11'd663: sine = 32'h3f650479;
    11'd664: sine = 32'h3f64aa59;
    11'd665: sine = 32'h3f644fac;
    11'd666: sine = 32'h3f63f473;
    11'd667: sine = 32'h3f6398ad;
    11'd668: sine = 32'h3f633c5a;
    11'd669: sine = 32'h3f62df7b;
    11'd670: sine = 32'h3f628210;
    11'd671: sine = 32'h3f62241a;
    11'd672: sine = 32'h3f61c598;
    11'd673: sine = 32'h3f61668b;
    11'd674: sine = 32'h3f6106f2;
    11'd675: sine = 32'h3f60a6cf;
    11'd676: sine = 32'h3f604621;
    11'd677: sine = 32'h3f5fe4e9;
    11'd678: sine = 32'h3f5f8327;
    11'd679: sine = 32'h3f5f20db;
    11'd680: sine = 32'h3f5ebe06;
    11'd681: sine = 32'h3f5e5aa7;
    11'd682: sine = 32'h3f5df6be;
    11'd683: sine = 32'h3f5d924d;
    11'd684: sine = 32'h3f5d2d54;
    11'd685: sine = 32'h3f5cc7d1;
    11'd686: sine = 32'h3f5c61c7;
    11'd687: sine = 32'h3f5bfb35;
    11'd688: sine = 32'h3f5b941a;
    11'd689: sine = 32'h3f5b2c79;
    11'd690: sine = 32'h3f5ac450;
    11'd691: sine = 32'h3f5a5ba1;
    11'd692: sine = 32'h3f59f26a;
    11'd693: sine = 32'h3f5988ae;
    11'd694: sine = 32'h3f591e6b;
    11'd695: sine = 32'h3f58b3a2;
    11'd696: sine = 32'h3f584853;
    11'd697: sine = 32'h3f57dc7f;
    11'd698: sine = 32'h3f577026;
    11'd699: sine = 32'h3f570348;
    11'd700: sine = 32'h3f5695e5;
    11'd701: sine = 32'h3f5627fe;
    11'd702: sine = 32'h3f55b993;
    11'd703: sine = 32'h3f554aa4;
    11'd704: sine = 32'h3f54db32;
    11'd705: sine = 32'h3f546b3c;
    11'd706: sine = 32'h3f53fac3;
    11'd707: sine = 32'h3f5389c7;
    11'd708: sine = 32'h3f531849;
    11'd709: sine = 32'h3f52a649;
    11'd710: sine = 32'h3f5233c7;
    11'd711: sine = 32'h3f51c0c3;
    11'd712: sine = 32'h3f514d3d;
    11'd713: sine = 32'h3f50d937;
    11'd714: sine = 32'h3f5064b0;
    11'd715: sine = 32'h3f4fefa8;
    11'd716: sine = 32'h3f4f7a20;
    11'd717: sine = 32'h3f4f0418;
    11'd718: sine = 32'h3f4e8d90;
    11'd719: sine = 32'h3f4e1689;
    11'd720: sine = 32'h3f4d9f03;
    11'd721: sine = 32'h3f4d26fe;
    11'd722: sine = 32'h3f4cae7a;
    11'd723: sine = 32'h3f4c3578;
    11'd724: sine = 32'h3f4bbbf8;
    11'd725: sine = 32'h3f4b41fa;
    11'd726: sine = 32'h3f4ac780;
    11'd727: sine = 32'h3f4a4c88;
    11'd728: sine = 32'h3f49d113;
    11'd729: sine = 32'h3f495521;
    11'd730: sine = 32'h3f48d8b4;
    11'd731: sine = 32'h3f485bcb;
    11'd732: sine = 32'h3f47de66;
    11'd733: sine = 32'h3f476085;
    11'd734: sine = 32'h3f46e22a;
    11'd735: sine = 32'h3f466354;
    11'd736: sine = 32'h3f45e404;
    11'd737: sine = 32'h3f456439;
    11'd738: sine = 32'h3f44e3f5;
    11'd739: sine = 32'h3f446338;
    11'd740: sine = 32'h3f43e201;
    11'd741: sine = 32'h3f436051;
    11'd742: sine = 32'h3f42de29;
    11'd743: sine = 32'h3f425b89;
    11'd744: sine = 32'h3f41d871;
    11'd745: sine = 32'h3f4154e1;
    11'd746: sine = 32'h3f40d0da;
    11'd747: sine = 32'h3f404c5c;
    11'd748: sine = 32'h3f3fc768;
    11'd749: sine = 32'h3f3f41fd;
    11'd750: sine = 32'h3f3ebc1c;
    11'd751: sine = 32'h3f3e35c5;
    11'd752: sine = 32'h3f3daefa;
    11'd753: sine = 32'h3f3d27b9;
    11'd754: sine = 32'h3f3ca003;
    11'd755: sine = 32'h3f3c17d9;
    11'd756: sine = 32'h3f3b8f3b;
    11'd757: sine = 32'h3f3b062a;
    11'd758: sine = 32'h3f3a7ca5;
    11'd759: sine = 32'h3f39f2ad;
    11'd760: sine = 32'h3f396842;
    11'd761: sine = 32'h3f38dd65;
    11'd762: sine = 32'h3f385216;
    11'd763: sine = 32'h3f37c655;
    11'd764: sine = 32'h3f373a23;
    11'd765: sine = 32'h3f36ad80;
    11'd766: sine = 32'h3f36206c;
    11'd767: sine = 32'h3f3592e8;
    11'd768: sine = 32'h3f3504f4;
    11'd769: sine = 32'h3f347690;
    11'd770: sine = 32'h3f33e7bd;
    11'd771: sine = 32'h3f33587a;
    11'd772: sine = 32'h3f32c8ca;
    11'd773: sine = 32'h3f3238ab;
    11'd774: sine = 32'h3f31a81e;
    11'd775: sine = 32'h3f311723;
    11'd776: sine = 32'h3f3085bb;
    11'd777: sine = 32'h3f2ff3e6;
    11'd778: sine = 32'h3f2f61a5;
    11'd779: sine = 32'h3f2ecef8;
    11'd780: sine = 32'h3f2e3bde;
    11'd781: sine = 32'h3f2da85a;
    11'd782: sine = 32'h3f2d146a;
    11'd783: sine = 32'h3f2c800f;
    11'd784: sine = 32'h3f2beb4a;
    11'd785: sine = 32'h3f2b561b;
    11'd786: sine = 32'h3f2ac082;
    11'd787: sine = 32'h3f2a2a80;
    11'd788: sine = 32'h3f299415;
    11'd789: sine = 32'h3f28fd41;
    11'd790: sine = 32'h3f286606;
    11'd791: sine = 32'h3f27ce62;
    11'd792: sine = 32'h3f273656;
    11'd793: sine = 32'h3f269de4;
    11'd794: sine = 32'h3f26050b;
    11'd795: sine = 32'h3f256bcb;
    11'd796: sine = 32'h3f24d225;
    11'd797: sine = 32'h3f24381a;
    11'd798: sine = 32'h3f239da9;
    11'd799: sine = 32'h3f2302d4;
    11'd800: sine = 32'h3f22679a;
    11'd801: sine = 32'h3f21cbfb;
    11'd802: sine = 32'h3f212ff9;
    11'd803: sine = 32'h3f209394;
    11'd804: sine = 32'h3f1ff6cb;
    11'd805: sine = 32'h3f1f59a0;
    11'd806: sine = 32'h3f1ebc12;
    11'd807: sine = 32'h3f1e1e23;
    11'd808: sine = 32'h3f1d7fd2;
    11'd809: sine = 32'h3f1ce120;
    11'd810: sine = 32'h3f1c420d;
    11'd811: sine = 32'h3f1ba299;
    11'd812: sine = 32'h3f1b02c6;
    11'd813: sine = 32'h3f1a6293;
    11'd814: sine = 32'h3f19c201;
    11'd815: sine = 32'h3f192110;
    11'd816: sine = 32'h3f187fc0;
    11'd817: sine = 32'h3f17de13;
    11'd818: sine = 32'h3f173c08;
    11'd819: sine = 32'h3f16999f;
    11'd820: sine = 32'h3f15f6da;
    11'd821: sine = 32'h3f1553b8;
    11'd822: sine = 32'h3f14b03a;
    11'd823: sine = 32'h3f140c60;
    11'd824: sine = 32'h3f13682b;
    11'd825: sine = 32'h3f12c39b;
    11'd826: sine = 32'h3f121eb0;
    11'd827: sine = 32'h3f11796c;
    11'd828: sine = 32'h3f10d3cd;
    11'd829: sine = 32'h3f102dd6;
    11'd830: sine = 32'h3f0f8785;
    11'd831: sine = 32'h3f0ee0dc;
    11'd832: sine = 32'h3f0e39da;
    11'd833: sine = 32'h3f0d9281;
    11'd834: sine = 32'h3f0cead1;
    11'd835: sine = 32'h3f0c42ca;
    11'd836: sine = 32'h3f0b9a6c;
    11'd837: sine = 32'h3f0af1b8;
    11'd838: sine = 32'h3f0a48ae;
    11'd839: sine = 32'h3f099f4f;
    11'd840: sine = 32'h3f08f59b;
    11'd841: sine = 32'h3f084b93;
    11'd842: sine = 32'h3f07a136;
    11'd843: sine = 32'h3f06f686;
    11'd844: sine = 32'h3f064b83;
    11'd845: sine = 32'h3f05a02d;
    11'd846: sine = 32'h3f04f484;
    11'd847: sine = 32'h3f04488a;
    11'd848: sine = 32'h3f039c3d;
    11'd849: sine = 32'h3f02efa0;
    11'd850: sine = 32'h3f0242b2;
    11'd851: sine = 32'h3f019573;
    11'd852: sine = 32'h3f00e7e5;
    11'd853: sine = 32'h3f003a07;
    11'd854: sine = 32'h3eff17b4;
    11'd855: sine = 32'h3efdbabc;
    11'd856: sine = 32'h3efc5d28;
    11'd857: sine = 32'h3efafef9;
    11'd858: sine = 32'h3ef9a02e;
    11'd859: sine = 32'h3ef840ca;
    11'd860: sine = 32'h3ef6e0cc;
    11'd861: sine = 32'h3ef58036;
    11'd862: sine = 32'h3ef41f09;
    11'd863: sine = 32'h3ef2bd45;
    11'd864: sine = 32'h3ef15aeb;
    11'd865: sine = 32'h3eeff7fd;
    11'd866: sine = 32'h3eee947a;
    11'd867: sine = 32'h3eed3064;
    11'd868: sine = 32'h3eebcbbc;
    11'd869: sine = 32'h3eea6683;
    11'd870: sine = 32'h3ee900b9;
    11'd871: sine = 32'h3ee79a5f;
    11'd872: sine = 32'h3ee63376;
    11'd873: sine = 32'h3ee4cbff;
    11'd874: sine = 32'h3ee363fc;
    11'd875: sine = 32'h3ee1fb6c;
    11'd876: sine = 32'h3ee09250;
    11'd877: sine = 32'h3edf28aa;
    11'd878: sine = 32'h3eddbe7a;
    11'd879: sine = 32'h3edc53c2;
    11'd880: sine = 32'h3edae882;
    11'd881: sine = 32'h3ed97cba;
    11'd882: sine = 32'h3ed8106d;
    11'd883: sine = 32'h3ed6a39a;
    11'd884: sine = 32'h3ed53643;
    11'd885: sine = 32'h3ed3c868;
    11'd886: sine = 32'h3ed25a0b;
    11'd887: sine = 32'h3ed0eb2c;
    11'd888: sine = 32'h3ecf7bcc;
    11'd889: sine = 32'h3ece0bec;
    11'd890: sine = 32'h3ecc9b8c;
    11'd891: sine = 32'h3ecb2aaf;
    11'd892: sine = 32'h3ec9b955;
    11'd893: sine = 32'h3ec8477e;
    11'd894: sine = 32'h3ec6d52b;
    11'd895: sine = 32'h3ec5625e;
    11'd896: sine = 32'h3ec3ef17;
    11'd897: sine = 32'h3ec27b57;
    11'd898: sine = 32'h3ec1071f;
    11'd899: sine = 32'h3ebf9270;
    11'd900: sine = 32'h3ebe1d4b;
    11'd901: sine = 32'h3ebca7b1;
    11'd902: sine = 32'h3ebb31a2;
    11'd903: sine = 32'h3eb9bb20;
    11'd904: sine = 32'h3eb8442b;
    11'd905: sine = 32'h3eb6ccc5;
    11'd906: sine = 32'h3eb554ed;
    11'd907: sine = 32'h3eb3dca6;
    11'd908: sine = 32'h3eb263f0;
    11'd909: sine = 32'h3eb0eacc;
    11'd910: sine = 32'h3eaf713b;
    11'd911: sine = 32'h3eadf73e;
    11'd912: sine = 32'h3eac7cd5;
    11'd913: sine = 32'h3eab0202;
    11'd914: sine = 32'h3ea986c6;
    11'd915: sine = 32'h3ea80b20;
    11'd916: sine = 32'h3ea68f14;
    11'd917: sine = 32'h3ea512a0;
    11'd918: sine = 32'h3ea395c7;
    11'd919: sine = 32'h3ea21888;
    11'd920: sine = 32'h3ea09ae6;
    11'd921: sine = 32'h3e9f1ce1;
    11'd922: sine = 32'h3e9d9e79;
    11'd923: sine = 32'h3e9c1fb1;
    11'd924: sine = 32'h3e9aa088;
    11'd925: sine = 32'h3e9920ff;
    11'd926: sine = 32'h3e97a118;
    11'd927: sine = 32'h3e9620d4;
    11'd928: sine = 32'h3e94a033;
    11'd929: sine = 32'h3e931f36;
    11'd930: sine = 32'h3e919ddf;
    11'd931: sine = 32'h3e901c2e;
    11'd932: sine = 32'h3e8e9a24;
    11'd933: sine = 32'h3e8d17c1;
    11'd934: sine = 32'h3e8b9508;
    11'd935: sine = 32'h3e8a11f9;
    11'd936: sine = 32'h3e888e95;
    11'd937: sine = 32'h3e870adc;
    11'd938: sine = 32'h3e8586d0;
    11'd939: sine = 32'h3e840272;
    11'd940: sine = 32'h3e827dc2;
    11'd941: sine = 32'h3e80f8c2;
    11'd942: sine = 32'h3e7ee6e4;
    11'd943: sine = 32'h3e7bdba7;
    11'd944: sine = 32'h3e78cfcf;
    11'd945: sine = 32'h3e75c35d;
    11'd946: sine = 32'h3e72b654;
    11'd947: sine = 32'h3e6fa8b5;
    11'd948: sine = 32'h3e6c9a82;
    11'd949: sine = 32'h3e698bbe;
    11'd950: sine = 32'h3e667c69;
    11'd951: sine = 32'h3e636c86;
    11'd952: sine = 32'h3e605c17;
    11'd953: sine = 32'h3e5d4b1d;
    11'd954: sine = 32'h3e5a399b;
    11'd955: sine = 32'h3e572792;
    11'd956: sine = 32'h3e541504;
    11'd957: sine = 32'h3e5101f4;
    11'd958: sine = 32'h3e4dee63;
    11'd959: sine = 32'h3e4ada53;
    11'd960: sine = 32'h3e47c5c5;
    11'd961: sine = 32'h3e44b0bd;
    11'd962: sine = 32'h3e419b3b;
    11'd963: sine = 32'h3e3e8541;
    11'd964: sine = 32'h3e3b6ed2;
    11'd965: sine = 32'h3e3857f0;
    11'd966: sine = 32'h3e35409b;
    11'd967: sine = 32'h3e3228d7;
    11'd968: sine = 32'h3e2f10a5;
    11'd969: sine = 32'h3e2bf808;
    11'd970: sine = 32'h3e28df00;
    11'd971: sine = 32'h3e25c58f;
    11'd972: sine = 32'h3e22abb9;
    11'd973: sine = 32'h3e1f917e;
    11'd974: sine = 32'h3e1c76e1;
    11'd975: sine = 32'h3e195be3;
    11'd976: sine = 32'h3e164087;
    11'd977: sine = 32'h3e1324ce;
    11'd978: sine = 32'h3e1008ba;
    11'd979: sine = 32'h3e0cec4d;
    11'd980: sine = 32'h3e09cf8a;
    11'd981: sine = 32'h3e06b271;
    11'd982: sine = 32'h3e039506;
    11'd983: sine = 32'h3e007749;
    11'd984: sine = 32'h3dfab27a;
    11'd985: sine = 32'h3df475c7;
    11'd986: sine = 32'h3dee387d;
    11'd987: sine = 32'h3de7faa1;
    11'd988: sine = 32'h3de1bc35;
    11'd989: sine = 32'h3ddb7d3e;
    11'd990: sine = 32'h3dd53dc0;
    11'd991: sine = 32'h3dcefdbe;
    11'd992: sine = 32'h3dc8bd3d;
    11'd993: sine = 32'h3dc27c40;
    11'd994: sine = 32'h3dbc3aca;
    11'd995: sine = 32'h3db5f8e1;
    11'd996: sine = 32'h3dafb687;
    11'd997: sine = 32'h3da973c1;
    11'd998: sine = 32'h3da33093;
    11'd999: sine = 32'h3d9ced00;
    11'd1000: sine = 32'h3d96a90c;
    11'd1001: sine = 32'h3d9064bb;
    11'd1002: sine = 32'h3d8a2011;
    11'd1003: sine = 32'h3d83db11;
    11'd1004: sine = 32'h3d7b2b82;
    11'd1005: sine = 32'h3d6ea046;
    11'd1006: sine = 32'h3d621477;
    11'd1007: sine = 32'h3d55881c;
    11'd1008: sine = 32'h3d48fb3e;
    11'd1009: sine = 32'h3d3c6de3;
    11'd1010: sine = 32'h3d2fe015;
    11'd1011: sine = 32'h3d2351da;
    11'd1012: sine = 32'h3d16c33a;
    11'd1013: sine = 32'h3d0a343d;
    11'd1014: sine = 32'h3cfb49d6;
    11'd1015: sine = 32'h3ce22a97;
    11'd1016: sine = 32'h3cc90acc;
    11'd1017: sine = 32'h3cafea86;
    11'd1018: sine = 32'h3c96c9d2;
    11'd1019: sine = 32'h3c7b5185;
    11'd1020: sine = 32'h3c490ec9;
    11'd1021: sine = 32'h3c16cb92;
    11'd1022: sine = 32'h3bc90ffb;
    11'd1023: sine = 32'h3b4910ac;
    11'd1024: sine = 32'h33662a9a;
    11'd1025: sine = 32'hbb490ee0;
    11'd1026: sine = 32'hbbc90f15;
    11'd1027: sine = 32'hbc16cb1f;
    11'd1028: sine = 32'hbc490e56;
    11'd1029: sine = 32'hbc7b5112;
    11'd1030: sine = 32'hbc96c999;
    11'd1031: sine = 32'hbcafea4c;
    11'd1032: sine = 32'hbcc90a93;
    11'd1033: sine = 32'hbce22a5d;
    11'd1034: sine = 32'hbcfb499d;
    11'd1035: sine = 32'hbd0a3420;
    11'd1036: sine = 32'hbd16c31d;
    11'd1037: sine = 32'hbd2351bd;
    11'd1038: sine = 32'hbd2fdff8;
    11'd1039: sine = 32'hbd3c6dc7;
    11'd1040: sine = 32'hbd48fb21;
    11'd1041: sine = 32'hbd5587ff;
    11'd1042: sine = 32'hbd62145a;
    11'd1043: sine = 32'hbd6ea029;
    11'd1044: sine = 32'hbd7b2b65;
    11'd1045: sine = 32'hbd83db03;
    11'd1046: sine = 32'hbd8a2002;
    11'd1047: sine = 32'hbd9064ac;
    11'd1048: sine = 32'hbd96a8fd;
    11'd1049: sine = 32'hbd9cecf1;
    11'd1050: sine = 32'hbda33084;
    11'd1051: sine = 32'hbda973b3;
    11'd1052: sine = 32'hbdafb679;
    11'd1053: sine = 32'hbdb5f8d3;
    11'd1054: sine = 32'hbdbc3abc;
    11'd1055: sine = 32'hbdc27c31;
    11'd1056: sine = 32'hbdc8bd2e;
    11'd1057: sine = 32'hbdcefdb0;
    11'd1058: sine = 32'hbdd53db2;
    11'd1059: sine = 32'hbddb7d30;
    11'd1060: sine = 32'hbde1bc27;
    11'd1061: sine = 32'hbde7fa92;
    11'd1062: sine = 32'hbdee386f;
    11'd1063: sine = 32'hbdf475b9;
    11'd1064: sine = 32'hbdfab26b;
    11'd1065: sine = 32'hbe007742;
    11'd1066: sine = 32'hbe0394ff;
    11'd1067: sine = 32'hbe06b26a;
    11'd1068: sine = 32'hbe09cf83;
    11'd1069: sine = 32'hbe0cec46;
    11'd1070: sine = 32'hbe1008b3;
    11'd1071: sine = 32'hbe1324c7;
    11'd1072: sine = 32'hbe164080;
    11'd1073: sine = 32'hbe195bdc;
    11'd1074: sine = 32'hbe1c76da;
    11'd1075: sine = 32'hbe1f9177;
    11'd1076: sine = 32'hbe22abb2;
    11'd1077: sine = 32'hbe25c588;
    11'd1078: sine = 32'hbe28def8;
    11'd1079: sine = 32'hbe2bf800;
    11'd1080: sine = 32'hbe2f109e;
    11'd1081: sine = 32'hbe3228d0;
    11'd1082: sine = 32'hbe354094;
    11'd1083: sine = 32'hbe3857e9;
    11'd1084: sine = 32'hbe3b6ecb;
    11'd1085: sine = 32'hbe3e853a;
    11'd1086: sine = 32'hbe419b34;
    11'd1087: sine = 32'hbe44b0b5;
    11'd1088: sine = 32'hbe47c5be;
    11'd1089: sine = 32'hbe4ada4c;
    11'd1090: sine = 32'hbe4dee5c;
    11'd1091: sine = 32'hbe5101ed;
    11'd1092: sine = 32'hbe5414fd;
    11'd1093: sine = 32'hbe57278b;
    11'd1094: sine = 32'hbe5a3994;
    11'd1095: sine = 32'hbe5d4b16;
    11'd1096: sine = 32'hbe605c10;
    11'd1097: sine = 32'hbe636c7f;
    11'd1098: sine = 32'hbe667c62;
    11'd1099: sine = 32'hbe698bb7;
    11'd1100: sine = 32'hbe6c9a7b;
    11'd1101: sine = 32'hbe6fa8ae;
    11'd1102: sine = 32'hbe72b64d;
    11'd1103: sine = 32'hbe75c356;
    11'd1104: sine = 32'hbe78cfc8;
    11'd1105: sine = 32'hbe7bdba0;
    11'd1106: sine = 32'hbe7ee6dd;
    11'd1107: sine = 32'hbe80f8be;
    11'd1108: sine = 32'hbe827dbf;
    11'd1109: sine = 32'hbe84026e;
    11'd1110: sine = 32'hbe8586cd;
    11'd1111: sine = 32'hbe870ad9;
    11'd1112: sine = 32'hbe888e91;
    11'd1113: sine = 32'hbe8a11f6;
    11'd1114: sine = 32'hbe8b9505;
    11'd1115: sine = 32'hbe8d17be;
    11'd1116: sine = 32'hbe8e9a20;
    11'd1117: sine = 32'hbe901c2a;
    11'd1118: sine = 32'hbe919ddb;
    11'd1119: sine = 32'hbe931f33;
    11'd1120: sine = 32'hbe94a030;
    11'd1121: sine = 32'hbe9620d1;
    11'd1122: sine = 32'hbe97a115;
    11'd1123: sine = 32'hbe9920fc;
    11'd1124: sine = 32'hbe9aa084;
    11'd1125: sine = 32'hbe9c1fad;
    11'd1126: sine = 32'hbe9d9e76;
    11'd1127: sine = 32'hbe9f1cdd;
    11'd1128: sine = 32'hbea09ae3;
    11'd1129: sine = 32'hbea21885;
    11'd1130: sine = 32'hbea395c3;
    11'd1131: sine = 32'hbea5129d;
    11'd1132: sine = 32'hbea68f10;
    11'd1133: sine = 32'hbea80b1d;
    11'd1134: sine = 32'hbea986c2;
    11'd1135: sine = 32'hbeab01ff;
    11'd1136: sine = 32'hbeac7cd2;
    11'd1137: sine = 32'hbeadf73a;
    11'd1138: sine = 32'hbeaf7138;
    11'd1139: sine = 32'hbeb0eac9;
    11'd1140: sine = 32'hbeb263ed;
    11'd1141: sine = 32'hbeb3dca3;
    11'd1142: sine = 32'hbeb554ea;
    11'd1143: sine = 32'hbeb6ccc1;
    11'd1144: sine = 32'hbeb84428;
    11'd1145: sine = 32'hbeb9bb1c;
    11'd1146: sine = 32'hbebb319f;
    11'd1147: sine = 32'hbebca7ad;
    11'd1148: sine = 32'hbebe1d48;
    11'd1149: sine = 32'hbebf926d;
    11'd1150: sine = 32'hbec1071c;
    11'd1151: sine = 32'hbec27b53;
    11'd1152: sine = 32'hbec3ef13;
    11'd1153: sine = 32'hbec5625a;
    11'd1154: sine = 32'hbec6d528;
    11'd1155: sine = 32'hbec8477a;
    11'd1156: sine = 32'hbec9b951;
    11'd1157: sine = 32'hbecb2aac;
    11'd1158: sine = 32'hbecc9b89;
    11'd1159: sine = 32'hbece0be8;
    11'd1160: sine = 32'hbecf7bc8;
    11'd1161: sine = 32'hbed0eb28;
    11'd1162: sine = 32'hbed25a07;
    11'd1163: sine = 32'hbed3c865;
    11'd1164: sine = 32'hbed5363f;
    11'd1165: sine = 32'hbed6a397;
    11'd1166: sine = 32'hbed8106a;
    11'd1167: sine = 32'hbed97cb7;
    11'd1168: sine = 32'hbedae87e;
    11'd1169: sine = 32'hbedc53bf;
    11'd1170: sine = 32'hbeddbe77;
    11'd1171: sine = 32'hbedf28a7;
    11'd1172: sine = 32'hbee0924d;
    11'd1173: sine = 32'hbee1fb68;
    11'd1174: sine = 32'hbee363f8;
    11'd1175: sine = 32'hbee4cbfc;
    11'd1176: sine = 32'hbee63373;
    11'd1177: sine = 32'hbee79a5c;
    11'd1178: sine = 32'hbee900b5;
    11'd1179: sine = 32'hbeea6680;
    11'd1180: sine = 32'hbeebcbb9;
    11'd1181: sine = 32'hbeed3061;
    11'd1182: sine = 32'hbeee9477;
    11'd1183: sine = 32'hbeeff7f9;
    11'd1184: sine = 32'hbef15ae8;
    11'd1185: sine = 32'hbef2bd42;
    11'd1186: sine = 32'hbef41f06;
    11'd1187: sine = 32'hbef58033;
    11'd1188: sine = 32'hbef6e0c9;
    11'd1189: sine = 32'hbef840c6;
    11'd1190: sine = 32'hbef9a02b;
    11'd1191: sine = 32'hbefafef5;
    11'd1192: sine = 32'hbefc5d25;
    11'd1193: sine = 32'hbefdbab9;
    11'd1194: sine = 32'hbeff17b1;
    11'd1195: sine = 32'hbf003a05;
    11'd1196: sine = 32'hbf00e7e3;
    11'd1197: sine = 32'hbf019572;
    11'd1198: sine = 32'hbf0242b0;
    11'd1199: sine = 32'hbf02ef9e;
    11'd1200: sine = 32'hbf039c3c;
    11'd1201: sine = 32'hbf044888;
    11'd1202: sine = 32'hbf04f483;
    11'd1203: sine = 32'hbf05a02b;
    11'd1204: sine = 32'hbf064b82;
    11'd1205: sine = 32'hbf06f685;
    11'd1206: sine = 32'hbf07a135;
    11'd1207: sine = 32'hbf084b91;
    11'd1208: sine = 32'hbf08f59a;
    11'd1209: sine = 32'hbf099f4e;
    11'd1210: sine = 32'hbf0a48ad;
    11'd1211: sine = 32'hbf0af1b6;
    11'd1212: sine = 32'hbf0b9a6a;
    11'd1213: sine = 32'hbf0c42c8;
    11'd1214: sine = 32'hbf0ceacf;
    11'd1215: sine = 32'hbf0d9280;
    11'd1216: sine = 32'hbf0e39d9;
    11'd1217: sine = 32'hbf0ee0da;
    11'd1218: sine = 32'hbf0f8783;
    11'd1219: sine = 32'hbf102dd4;
    11'd1220: sine = 32'hbf10d3cc;
    11'd1221: sine = 32'hbf11796a;
    11'd1222: sine = 32'hbf121eaf;
    11'd1223: sine = 32'hbf12c39a;
    11'd1224: sine = 32'hbf13682a;
    11'd1225: sine = 32'hbf140c5f;
    11'd1226: sine = 32'hbf14b038;
    11'd1227: sine = 32'hbf1553b6;
    11'd1228: sine = 32'hbf15f6d8;
    11'd1229: sine = 32'hbf16999e;
    11'd1230: sine = 32'hbf173c06;
    11'd1231: sine = 32'hbf17de11;
    11'd1232: sine = 32'hbf187fbf;
    11'd1233: sine = 32'hbf19210f;
    11'd1234: sine = 32'hbf19c200;
    11'd1235: sine = 32'hbf1a6292;
    11'd1236: sine = 32'hbf1b02c5;
    11'd1237: sine = 32'hbf1ba298;
    11'd1238: sine = 32'hbf1c420b;
    11'd1239: sine = 32'hbf1ce11e;
    11'd1240: sine = 32'hbf1d7fd0;
    11'd1241: sine = 32'hbf1e1e21;
    11'd1242: sine = 32'hbf1ebc11;
    11'd1243: sine = 32'hbf1f599e;
    11'd1244: sine = 32'hbf1ff6ca;
    11'd1245: sine = 32'hbf209392;
    11'd1246: sine = 32'hbf212ff8;
    11'd1247: sine = 32'hbf21cbfa;
    11'd1248: sine = 32'hbf226798;
    11'd1249: sine = 32'hbf2302d2;
    11'd1250: sine = 32'hbf239da8;
    11'd1251: sine = 32'hbf243819;
    11'd1252: sine = 32'hbf24d224;
    11'd1253: sine = 32'hbf256bca;
    11'd1254: sine = 32'hbf260509;
    11'd1255: sine = 32'hbf269de3;
    11'd1256: sine = 32'hbf273655;
    11'd1257: sine = 32'hbf27ce60;
    11'd1258: sine = 32'hbf286604;
    11'd1259: sine = 32'hbf28fd40;
    11'd1260: sine = 32'hbf299414;
    11'd1261: sine = 32'hbf2a2a7f;
    11'd1262: sine = 32'hbf2ac081;
    11'd1263: sine = 32'hbf2b561a;
    11'd1264: sine = 32'hbf2beb49;
    11'd1265: sine = 32'hbf2c800e;
    11'd1266: sine = 32'hbf2d1469;
    11'd1267: sine = 32'hbf2da858;
    11'd1268: sine = 32'hbf2e3bdd;
    11'd1269: sine = 32'hbf2ecef6;
    11'd1270: sine = 32'hbf2f61a4;
    11'd1271: sine = 32'hbf2ff3e5;
    11'd1272: sine = 32'hbf3085ba;
    11'd1273: sine = 32'hbf311722;
    11'd1274: sine = 32'hbf31a81c;
    11'd1275: sine = 32'hbf3238a9;
    11'd1276: sine = 32'hbf32c8c8;
    11'd1277: sine = 32'hbf335879;
    11'd1278: sine = 32'hbf33e7bb;
    11'd1279: sine = 32'hbf34768f;
    11'd1280: sine = 32'hbf3504f2;
    11'd1281: sine = 32'hbf3592e7;
    11'd1282: sine = 32'hbf36206b;
    11'd1283: sine = 32'hbf36ad7f;
    11'd1284: sine = 32'hbf373a22;
    11'd1285: sine = 32'hbf37c654;
    11'd1286: sine = 32'hbf385215;
    11'd1287: sine = 32'hbf38dd64;
    11'd1288: sine = 32'hbf396841;
    11'd1289: sine = 32'hbf39f2ac;
    11'd1290: sine = 32'hbf3a7ca4;
    11'd1291: sine = 32'hbf3b0629;
    11'd1292: sine = 32'hbf3b8f3a;
    11'd1293: sine = 32'hbf3c17d8;
    11'd1294: sine = 32'hbf3ca002;
    11'd1295: sine = 32'hbf3d27b7;
    11'd1296: sine = 32'hbf3daef8;
    11'd1297: sine = 32'hbf3e35c4;
    11'd1298: sine = 32'hbf3ebc1b;
    11'd1299: sine = 32'hbf3f41fb;
    11'd1300: sine = 32'hbf3fc766;
    11'd1301: sine = 32'hbf404c5b;
    11'd1302: sine = 32'hbf40d0d9;
    11'd1303: sine = 32'hbf4154e0;
    11'd1304: sine = 32'hbf41d870;
    11'd1305: sine = 32'hbf425b88;
    11'd1306: sine = 32'hbf42de28;
    11'd1307: sine = 32'hbf436050;
    11'd1308: sine = 32'hbf43e200;
    11'd1309: sine = 32'hbf446336;
    11'd1310: sine = 32'hbf44e3f4;
    11'd1311: sine = 32'hbf456438;
    11'd1312: sine = 32'hbf45e403;
    11'd1313: sine = 32'hbf466353;
    11'd1314: sine = 32'hbf46e229;
    11'd1315: sine = 32'hbf476084;
    11'd1316: sine = 32'hbf47de64;
    11'd1317: sine = 32'hbf485bc9;
    11'd1318: sine = 32'hbf48d8b3;
    11'd1319: sine = 32'hbf495520;
    11'd1320: sine = 32'hbf49d112;
    11'd1321: sine = 32'hbf4a4c86;
    11'd1322: sine = 32'hbf4ac77e;
    11'd1323: sine = 32'hbf4b41f9;
    11'd1324: sine = 32'hbf4bbbf7;
    11'd1325: sine = 32'hbf4c3577;
    11'd1326: sine = 32'hbf4cae79;
    11'd1327: sine = 32'hbf4d26fc;
    11'd1328: sine = 32'hbf4d9f02;
    11'd1329: sine = 32'hbf4e1688;
    11'd1330: sine = 32'hbf4e8d8f;
    11'd1331: sine = 32'hbf4f0417;
    11'd1332: sine = 32'hbf4f7a1f;
    11'd1333: sine = 32'hbf4fefa7;
    11'd1334: sine = 32'hbf5064af;
    11'd1335: sine = 32'hbf50d936;
    11'd1336: sine = 32'hbf514d3c;
    11'd1337: sine = 32'hbf51c0c2;
    11'd1338: sine = 32'hbf5233c6;
    11'd1339: sine = 32'hbf52a648;
    11'd1340: sine = 32'hbf531848;
    11'd1341: sine = 32'hbf5389c6;
    11'd1342: sine = 32'hbf53fac2;
    11'd1343: sine = 32'hbf546b3b;
    11'd1344: sine = 32'hbf54db31;
    11'd1345: sine = 32'hbf554aa3;
    11'd1346: sine = 32'hbf55b992;
    11'd1347: sine = 32'hbf5627fd;
    11'd1348: sine = 32'hbf5695e4;
    11'd1349: sine = 32'hbf570347;
    11'd1350: sine = 32'hbf577025;
    11'd1351: sine = 32'hbf57dc7e;
    11'd1352: sine = 32'hbf584852;
    11'd1353: sine = 32'hbf58b3a1;
    11'd1354: sine = 32'hbf591e6a;
    11'd1355: sine = 32'hbf5988ad;
    11'd1356: sine = 32'hbf59f269;
    11'd1357: sine = 32'hbf5a5ba0;
    11'd1358: sine = 32'hbf5ac44f;
    11'd1359: sine = 32'hbf5b2c78;
    11'd1360: sine = 32'hbf5b941a;
    11'd1361: sine = 32'hbf5bfb34;
    11'd1362: sine = 32'hbf5c61c6;
    11'd1363: sine = 32'hbf5cc7d0;
    11'd1364: sine = 32'hbf5d2d53;
    11'd1365: sine = 32'hbf5d924c;
    11'd1366: sine = 32'hbf5df6be;
    11'd1367: sine = 32'hbf5e5aa6;
    11'd1368: sine = 32'hbf5ebe05;
    11'd1369: sine = 32'hbf5f20da;
    11'd1370: sine = 32'hbf5f8326;
    11'd1371: sine = 32'hbf5fe4e9;
    11'd1372: sine = 32'hbf604621;
    11'd1373: sine = 32'hbf60a6ce;
    11'd1374: sine = 32'hbf6106f1;
    11'd1375: sine = 32'hbf61668a;
    11'd1376: sine = 32'hbf61c597;
    11'd1377: sine = 32'hbf622419;
    11'd1378: sine = 32'hbf62820f;
    11'd1379: sine = 32'hbf62df7a;
    11'd1380: sine = 32'hbf633c59;
    11'd1381: sine = 32'hbf6398ac;
    11'd1382: sine = 32'hbf63f472;
    11'd1383: sine = 32'hbf644fac;
    11'd1384: sine = 32'hbf64aa58;
    11'd1385: sine = 32'hbf650478;
    11'd1386: sine = 32'hbf655e0b;
    11'd1387: sine = 32'hbf65b710;
    11'd1388: sine = 32'hbf660f87;
    11'd1389: sine = 32'hbf666770;
    11'd1390: sine = 32'hbf66becc;
    11'd1391: sine = 32'hbf671599;
    11'd1392: sine = 32'hbf676bd7;
    11'd1393: sine = 32'hbf67c187;
    11'd1394: sine = 32'hbf6816a7;
    11'd1395: sine = 32'hbf686b39;
    11'd1396: sine = 32'hbf68bf3b;
    11'd1397: sine = 32'hbf6912ae;
    11'd1398: sine = 32'hbf696591;
    11'd1399: sine = 32'hbf69b7e3;
    11'd1400: sine = 32'hbf6a09a6;
    11'd1401: sine = 32'hbf6a5ad8;
    11'd1402: sine = 32'hbf6aab7a;
    11'd1403: sine = 32'hbf6afb8b;
    11'd1404: sine = 32'hbf6b4b0b;
    11'd1405: sine = 32'hbf6b99fa;
    11'd1406: sine = 32'hbf6be858;
    11'd1407: sine = 32'hbf6c3624;
    11'd1408: sine = 32'hbf6c835e;
    11'd1409: sine = 32'hbf6cd006;
    11'd1410: sine = 32'hbf6d1c1d;
    11'd1411: sine = 32'hbf6d67a1;
    11'd1412: sine = 32'hbf6db293;
    11'd1413: sine = 32'hbf6dfcf2;
    11'd1414: sine = 32'hbf6e46be;
    11'd1415: sine = 32'hbf6e8ff7;
    11'd1416: sine = 32'hbf6ed89d;
    11'd1417: sine = 32'hbf6f20b0;
    11'd1418: sine = 32'hbf6f682f;
    11'd1419: sine = 32'hbf6faf1b;
    11'd1420: sine = 32'hbf6ff573;
    11'd1421: sine = 32'hbf703b36;
    11'd1422: sine = 32'hbf708066;
    11'd1423: sine = 32'hbf70c501;
    11'd1424: sine = 32'hbf710908;
    11'd1425: sine = 32'hbf714c7a;
    11'd1426: sine = 32'hbf718f57;
    11'd1427: sine = 32'hbf71d19f;
    11'd1428: sine = 32'hbf721352;
    11'd1429: sine = 32'hbf725470;
    11'd1430: sine = 32'hbf7294f8;
    11'd1431: sine = 32'hbf72d4ea;
    11'd1432: sine = 32'hbf731447;
    11'd1433: sine = 32'hbf73530e;
    11'd1434: sine = 32'hbf73913e;
    11'd1435: sine = 32'hbf73ced9;
    11'd1436: sine = 32'hbf740bdd;
    11'd1437: sine = 32'hbf74484a;
    11'd1438: sine = 32'hbf748421;
    11'd1439: sine = 32'hbf74bf61;
    11'd1440: sine = 32'hbf74fa0a;
    11'd1441: sine = 32'hbf75341c;
    11'd1442: sine = 32'hbf756d97;
    11'd1443: sine = 32'hbf75a67a;
    11'd1444: sine = 32'hbf75dec6;
    11'd1445: sine = 32'hbf76167a;
    11'd1446: sine = 32'hbf764d96;
    11'd1447: sine = 32'hbf76841b;
    11'd1448: sine = 32'hbf76ba07;
    11'd1449: sine = 32'hbf76ef5b;
    11'd1450: sine = 32'hbf772417;
    11'd1451: sine = 32'hbf77583a;
    11'd1452: sine = 32'hbf778bc5;
    11'd1453: sine = 32'hbf77beb7;
    11'd1454: sine = 32'hbf77f110;
    11'd1455: sine = 32'hbf7822d0;
    11'd1456: sine = 32'hbf7853f8;
    11'd1457: sine = 32'hbf788486;
    11'd1458: sine = 32'hbf78b47a;
    11'd1459: sine = 32'hbf78e3d6;
    11'd1460: sine = 32'hbf791297;
    11'd1461: sine = 32'hbf7940c0;
    11'd1462: sine = 32'hbf796e4e;
    11'd1463: sine = 32'hbf799b43;
    11'd1464: sine = 32'hbf79c79d;
    11'd1465: sine = 32'hbf79f35e;
    11'd1466: sine = 32'hbf7a1e84;
    11'd1467: sine = 32'hbf7a4910;
    11'd1468: sine = 32'hbf7a7302;
    11'd1469: sine = 32'hbf7a9c59;
    11'd1470: sine = 32'hbf7ac515;
    11'd1471: sine = 32'hbf7aed37;
    11'd1472: sine = 32'hbf7b14be;
    11'd1473: sine = 32'hbf7b3baa;
    11'd1474: sine = 32'hbf7b61fc;
    11'd1475: sine = 32'hbf7b87b2;
    11'd1476: sine = 32'hbf7baccd;
    11'd1477: sine = 32'hbf7bd14d;
    11'd1478: sine = 32'hbf7bf531;
    11'd1479: sine = 32'hbf7c187a;
    11'd1480: sine = 32'hbf7c3b28;
    11'd1481: sine = 32'hbf7c5d3a;
    11'd1482: sine = 32'hbf7c7eb0;
    11'd1483: sine = 32'hbf7c9f8a;
    11'd1484: sine = 32'hbf7cbfc9;
    11'd1485: sine = 32'hbf7cdf6c;
    11'd1486: sine = 32'hbf7cfe72;
    11'd1487: sine = 32'hbf7d1cdd;
    11'd1488: sine = 32'hbf7d3aac;
    11'd1489: sine = 32'hbf7d57de;
    11'd1490: sine = 32'hbf7d7474;
    11'd1491: sine = 32'hbf7d906e;
    11'd1492: sine = 32'hbf7dabcb;
    11'd1493: sine = 32'hbf7dc68c;
    11'd1494: sine = 32'hbf7de0b1;
    11'd1495: sine = 32'hbf7dfa38;
    11'd1496: sine = 32'hbf7e1323;
    11'd1497: sine = 32'hbf7e2b72;
    11'd1498: sine = 32'hbf7e4323;
    11'd1499: sine = 32'hbf7e5a38;
    11'd1500: sine = 32'hbf7e70b0;
    11'd1501: sine = 32'hbf7e868b;
    11'd1502: sine = 32'hbf7e9bc8;
    11'd1503: sine = 32'hbf7eb069;
    11'd1504: sine = 32'hbf7ec46d;
    11'd1505: sine = 32'hbf7ed7d4;
    11'd1506: sine = 32'hbf7eea9d;
    11'd1507: sine = 32'hbf7efcc9;
    11'd1508: sine = 32'hbf7f0e58;
    11'd1509: sine = 32'hbf7f1f49;
    11'd1510: sine = 32'hbf7f2f9d;
    11'd1511: sine = 32'hbf7f3f54;
    11'd1512: sine = 32'hbf7f4e6d;
    11'd1513: sine = 32'hbf7f5ce9;
    11'd1514: sine = 32'hbf7f6ac7;
    11'd1515: sine = 32'hbf7f7808;
    11'd1516: sine = 32'hbf7f84ab;
    11'd1517: sine = 32'hbf7f90b1;
    11'd1518: sine = 32'hbf7f9c18;
    11'd1519: sine = 32'hbf7fa6e3;
    11'd1520: sine = 32'hbf7fb10f;
    11'd1521: sine = 32'hbf7fba9e;
    11'd1522: sine = 32'hbf7fc38f;
    11'd1523: sine = 32'hbf7fcbe2;
    11'd1524: sine = 32'hbf7fd397;
    11'd1525: sine = 32'hbf7fdaaf;
    11'd1526: sine = 32'hbf7fe129;
    11'd1527: sine = 32'hbf7fe705;
    11'd1528: sine = 32'hbf7fec43;
    11'd1529: sine = 32'hbf7ff0e3;
    11'd1530: sine = 32'hbf7ff4e6;
    11'd1531: sine = 32'hbf7ff84a;
    11'd1532: sine = 32'hbf7ffb11;
    11'd1533: sine = 32'hbf7ffd39;
    11'd1534: sine = 32'hbf7ffec4;
    11'd1535: sine = 32'hbf7fffb1;
    11'd1536: sine = 32'hbf800000;
    11'd1537: sine = 32'hbf7fffb1;
    11'd1538: sine = 32'hbf7ffec4;
    11'd1539: sine = 32'hbf7ffd39;
    11'd1540: sine = 32'hbf7ffb11;
    11'd1541: sine = 32'hbf7ff84a;
    11'd1542: sine = 32'hbf7ff4e6;
    11'd1543: sine = 32'hbf7ff0e3;
    11'd1544: sine = 32'hbf7fec43;
    11'd1545: sine = 32'hbf7fe705;
    11'd1546: sine = 32'hbf7fe129;
    11'd1547: sine = 32'hbf7fdaaf;
    11'd1548: sine = 32'hbf7fd398;
    11'd1549: sine = 32'hbf7fcbe2;
    11'd1550: sine = 32'hbf7fc38f;
    11'd1551: sine = 32'hbf7fba9e;
    11'd1552: sine = 32'hbf7fb10f;
    11'd1553: sine = 32'hbf7fa6e3;
    11'd1554: sine = 32'hbf7f9c19;
    11'd1555: sine = 32'hbf7f90b1;
    11'd1556: sine = 32'hbf7f84ab;
    11'd1557: sine = 32'hbf7f7808;
    11'd1558: sine = 32'hbf7f6ac7;
    11'd1559: sine = 32'hbf7f5ce9;
    11'd1560: sine = 32'hbf7f4e6e;
    11'd1561: sine = 32'hbf7f3f54;
    11'd1562: sine = 32'hbf7f2f9e;
    11'd1563: sine = 32'hbf7f1f49;
    11'd1564: sine = 32'hbf7f0e58;
    11'd1565: sine = 32'hbf7efcc9;
    11'd1566: sine = 32'hbf7eea9d;
    11'd1567: sine = 32'hbf7ed7d4;
    11'd1568: sine = 32'hbf7ec46d;
    11'd1569: sine = 32'hbf7eb06a;
    11'd1570: sine = 32'hbf7e9bc9;
    11'd1571: sine = 32'hbf7e868b;
    11'd1572: sine = 32'hbf7e70b0;
    11'd1573: sine = 32'hbf7e5a38;
    11'd1574: sine = 32'hbf7e4324;
    11'd1575: sine = 32'hbf7e2b72;
    11'd1576: sine = 32'hbf7e1324;
    11'd1577: sine = 32'hbf7dfa39;
    11'd1578: sine = 32'hbf7de0b1;
    11'd1579: sine = 32'hbf7dc68d;
    11'd1580: sine = 32'hbf7dabcc;
    11'd1581: sine = 32'hbf7d906e;
    11'd1582: sine = 32'hbf7d7475;
    11'd1583: sine = 32'hbf7d57df;
    11'd1584: sine = 32'hbf7d3aac;
    11'd1585: sine = 32'hbf7d1cde;
    11'd1586: sine = 32'hbf7cfe73;
    11'd1587: sine = 32'hbf7cdf6c;
    11'd1588: sine = 32'hbf7cbfc9;
    11'd1589: sine = 32'hbf7c9f8b;
    11'd1590: sine = 32'hbf7c7eb0;
    11'd1591: sine = 32'hbf7c5d3a;
    11'd1592: sine = 32'hbf7c3b28;
    11'd1593: sine = 32'hbf7c187b;
    11'd1594: sine = 32'hbf7bf532;
    11'd1595: sine = 32'hbf7bd14d;
    11'd1596: sine = 32'hbf7baccd;
    11'd1597: sine = 32'hbf7b87b2;
    11'd1598: sine = 32'hbf7b61fc;
    11'd1599: sine = 32'hbf7b3bab;
    11'd1600: sine = 32'hbf7b14bf;
    11'd1601: sine = 32'hbf7aed38;
    11'd1602: sine = 32'hbf7ac516;
    11'd1603: sine = 32'hbf7a9c59;
    11'd1604: sine = 32'hbf7a7302;
    11'd1605: sine = 32'hbf7a4911;
    11'd1606: sine = 32'hbf7a1e84;
    11'd1607: sine = 32'hbf79f35e;
    11'd1608: sine = 32'hbf79c79e;
    11'd1609: sine = 32'hbf799b43;
    11'd1610: sine = 32'hbf796e4f;
    11'd1611: sine = 32'hbf7940c0;
    11'd1612: sine = 32'hbf791298;
    11'd1613: sine = 32'hbf78e3d6;
    11'd1614: sine = 32'hbf78b47b;
    11'd1615: sine = 32'hbf788486;
    11'd1616: sine = 32'hbf7853f8;
    11'd1617: sine = 32'hbf7822d1;
    11'd1618: sine = 32'hbf77f111;
    11'd1619: sine = 32'hbf77beb8;
    11'd1620: sine = 32'hbf778bc5;
    11'd1621: sine = 32'hbf77583b;
    11'd1622: sine = 32'hbf772417;
    11'd1623: sine = 32'hbf76ef5c;
    11'd1624: sine = 32'hbf76ba08;
    11'd1625: sine = 32'hbf76841b;
    11'd1626: sine = 32'hbf764d97;
    11'd1627: sine = 32'hbf76167b;
    11'd1628: sine = 32'hbf75dec7;
    11'd1629: sine = 32'hbf75a67b;
    11'd1630: sine = 32'hbf756d98;
    11'd1631: sine = 32'hbf75341d;
    11'd1632: sine = 32'hbf74fa0b;
    11'd1633: sine = 32'hbf74bf62;
    11'd1634: sine = 32'hbf748422;
    11'd1635: sine = 32'hbf74484b;
    11'd1636: sine = 32'hbf740bde;
    11'd1637: sine = 32'hbf73ceda;
    11'd1638: sine = 32'hbf73913f;
    11'd1639: sine = 32'hbf73530f;
    11'd1640: sine = 32'hbf731448;
    11'd1641: sine = 32'hbf72d4eb;
    11'd1642: sine = 32'hbf7294f9;
    11'd1643: sine = 32'hbf725470;
    11'd1644: sine = 32'hbf721353;
    11'd1645: sine = 32'hbf71d1a0;
    11'd1646: sine = 32'hbf718f58;
    11'd1647: sine = 32'hbf714c7b;
    11'd1648: sine = 32'hbf710909;
    11'd1649: sine = 32'hbf70c502;
    11'd1650: sine = 32'hbf708067;
    11'd1651: sine = 32'hbf703b37;
    11'd1652: sine = 32'hbf6ff574;
    11'd1653: sine = 32'hbf6faf1c;
    11'd1654: sine = 32'hbf6f6830;
    11'd1655: sine = 32'hbf6f20b1;
    11'd1656: sine = 32'hbf6ed89e;
    11'd1657: sine = 32'hbf6e8ff8;
    11'd1658: sine = 32'hbf6e46bf;
    11'd1659: sine = 32'hbf6dfcf3;
    11'd1660: sine = 32'hbf6db294;
    11'd1661: sine = 32'hbf6d67a2;
    11'd1662: sine = 32'hbf6d1c1e;
    11'd1663: sine = 32'hbf6cd007;
    11'd1664: sine = 32'hbf6c835f;
    11'd1665: sine = 32'hbf6c3625;
    11'd1666: sine = 32'hbf6be859;
    11'd1667: sine = 32'hbf6b99fb;
    11'd1668: sine = 32'hbf6b4b0c;
    11'd1669: sine = 32'hbf6afb8c;
    11'd1670: sine = 32'hbf6aab7b;
    11'd1671: sine = 32'hbf6a5ad9;
    11'd1672: sine = 32'hbf6a09a7;
    11'd1673: sine = 32'hbf69b7e4;
    11'd1674: sine = 32'hbf696592;
    11'd1675: sine = 32'hbf6912af;
    11'd1676: sine = 32'hbf68bf3c;
    11'd1677: sine = 32'hbf686b3a;
    11'd1678: sine = 32'hbf6816a9;
    11'd1679: sine = 32'hbf67c188;
    11'd1680: sine = 32'hbf676bd8;
    11'd1681: sine = 32'hbf67159a;
    11'd1682: sine = 32'hbf66becd;
    11'd1683: sine = 32'hbf666772;
    11'd1684: sine = 32'hbf660f88;
    11'd1685: sine = 32'hbf65b711;
    11'd1686: sine = 32'hbf655e0c;
    11'd1687: sine = 32'hbf650479;
    11'd1688: sine = 32'hbf64aa5a;
    11'd1689: sine = 32'hbf644fad;
    11'd1690: sine = 32'hbf63f473;
    11'd1691: sine = 32'hbf6398ad;
    11'd1692: sine = 32'hbf633c5a;
    11'd1693: sine = 32'hbf62df7c;
    11'd1694: sine = 32'hbf628211;
    11'd1695: sine = 32'hbf62241a;
    11'd1696: sine = 32'hbf61c598;
    11'd1697: sine = 32'hbf61668b;
    11'd1698: sine = 32'hbf6106f3;
    11'd1699: sine = 32'hbf60a6d0;
    11'd1700: sine = 32'hbf604622;
    11'd1701: sine = 32'hbf5fe4ea;
    11'd1702: sine = 32'hbf5f8328;
    11'd1703: sine = 32'hbf5f20dc;
    11'd1704: sine = 32'hbf5ebe06;
    11'd1705: sine = 32'hbf5e5aa7;
    11'd1706: sine = 32'hbf5df6bf;
    11'd1707: sine = 32'hbf5d924e;
    11'd1708: sine = 32'hbf5d2d54;
    11'd1709: sine = 32'hbf5cc7d2;
    11'd1710: sine = 32'hbf5c61c7;
    11'd1711: sine = 32'hbf5bfb35;
    11'd1712: sine = 32'hbf5b941b;
    11'd1713: sine = 32'hbf5b2c79;
    11'd1714: sine = 32'hbf5ac451;
    11'd1715: sine = 32'hbf5a5ba1;
    11'd1716: sine = 32'hbf59f26b;
    11'd1717: sine = 32'hbf5988ae;
    11'd1718: sine = 32'hbf591e6b;
    11'd1719: sine = 32'hbf58b3a2;
    11'd1720: sine = 32'hbf584854;
    11'd1721: sine = 32'hbf57dc80;
    11'd1722: sine = 32'hbf577026;
    11'd1723: sine = 32'hbf570348;
    11'd1724: sine = 32'hbf5695e6;
    11'd1725: sine = 32'hbf5627ff;
    11'd1726: sine = 32'hbf55b994;
    11'd1727: sine = 32'hbf554aa5;
    11'd1728: sine = 32'hbf54db32;
    11'd1729: sine = 32'hbf546b3c;
    11'd1730: sine = 32'hbf53fac3;
    11'd1731: sine = 32'hbf5389c8;
    11'd1732: sine = 32'hbf53184a;
    11'd1733: sine = 32'hbf52a649;
    11'd1734: sine = 32'hbf5233c7;
    11'd1735: sine = 32'hbf51c0c3;
    11'd1736: sine = 32'hbf514d3e;
    11'd1737: sine = 32'hbf50d937;
    11'd1738: sine = 32'hbf5064b0;
    11'd1739: sine = 32'hbf4fefa8;
    11'd1740: sine = 32'hbf4f7a20;
    11'd1741: sine = 32'hbf4f0418;
    11'd1742: sine = 32'hbf4e8d91;
    11'd1743: sine = 32'hbf4e1689;
    11'd1744: sine = 32'hbf4d9f03;
    11'd1745: sine = 32'hbf4d26fe;
    11'd1746: sine = 32'hbf4cae7a;
    11'd1747: sine = 32'hbf4c3578;
    11'd1748: sine = 32'hbf4bbbf9;
    11'd1749: sine = 32'hbf4b41fb;
    11'd1750: sine = 32'hbf4ac780;
    11'd1751: sine = 32'hbf4a4c88;
    11'd1752: sine = 32'hbf49d113;
    11'd1753: sine = 32'hbf495522;
    11'd1754: sine = 32'hbf48d8b4;
    11'd1755: sine = 32'hbf485bcb;
    11'd1756: sine = 32'hbf47de66;
    11'd1757: sine = 32'hbf476086;
    11'd1758: sine = 32'hbf46e22b;
    11'd1759: sine = 32'hbf466355;
    11'd1760: sine = 32'hbf45e404;
    11'd1761: sine = 32'hbf45643a;
    11'd1762: sine = 32'hbf44e3f6;
    11'd1763: sine = 32'hbf446338;
    11'd1764: sine = 32'hbf43e201;
    11'd1765: sine = 32'hbf436052;
    11'd1766: sine = 32'hbf42de2a;
    11'd1767: sine = 32'hbf425b8a;
    11'd1768: sine = 32'hbf41d871;
    11'd1769: sine = 32'hbf4154e2;
    11'd1770: sine = 32'hbf40d0db;
    11'd1771: sine = 32'hbf404c5d;
    11'd1772: sine = 32'hbf3fc768;
    11'd1773: sine = 32'hbf3f41fd;
    11'd1774: sine = 32'hbf3ebc1c;
    11'd1775: sine = 32'hbf3e35c6;
    11'd1776: sine = 32'hbf3daefa;
    11'd1777: sine = 32'hbf3d27b9;
    11'd1778: sine = 32'hbf3ca004;
    11'd1779: sine = 32'hbf3c17da;
    11'd1780: sine = 32'hbf3b8f3c;
    11'd1781: sine = 32'hbf3b062a;
    11'd1782: sine = 32'hbf3a7ca5;
    11'd1783: sine = 32'hbf39f2ae;
    11'd1784: sine = 32'hbf396843;
    11'd1785: sine = 32'hbf38dd66;
    11'd1786: sine = 32'hbf385217;
    11'd1787: sine = 32'hbf37c656;
    11'd1788: sine = 32'hbf373a24;
    11'd1789: sine = 32'hbf36ad81;
    11'd1790: sine = 32'hbf36206d;
    11'd1791: sine = 32'hbf3592e9;
    11'd1792: sine = 32'hbf3504f4;
    11'd1793: sine = 32'hbf347690;
    11'd1794: sine = 32'hbf33e7bd;
    11'd1795: sine = 32'hbf33587b;
    11'd1796: sine = 32'hbf32c8ca;
    11'd1797: sine = 32'hbf3238ab;
    11'd1798: sine = 32'hbf31a81e;
    11'd1799: sine = 32'hbf311724;
    11'd1800: sine = 32'hbf3085bc;
    11'd1801: sine = 32'hbf2ff3e7;
    11'd1802: sine = 32'hbf2f61a6;
    11'd1803: sine = 32'hbf2ecef8;
    11'd1804: sine = 32'hbf2e3bdf;
    11'd1805: sine = 32'hbf2da85a;
    11'd1806: sine = 32'hbf2d146a;
    11'd1807: sine = 32'hbf2c8010;
    11'd1808: sine = 32'hbf2beb4b;
    11'd1809: sine = 32'hbf2b561c;
    11'd1810: sine = 32'hbf2ac083;
    11'd1811: sine = 32'hbf2a2a81;
    11'd1812: sine = 32'hbf299416;
    11'd1813: sine = 32'hbf28fd42;
    11'd1814: sine = 32'hbf286606;
    11'd1815: sine = 32'hbf27ce62;
    11'd1816: sine = 32'hbf273657;
    11'd1817: sine = 32'hbf269de5;
    11'd1818: sine = 32'hbf26050b;
    11'd1819: sine = 32'hbf256bcc;
    11'd1820: sine = 32'hbf24d226;
    11'd1821: sine = 32'hbf24381b;
    11'd1822: sine = 32'hbf239daa;
    11'd1823: sine = 32'hbf2302d5;
    11'd1824: sine = 32'hbf22679a;
    11'd1825: sine = 32'hbf21cbfc;
    11'd1826: sine = 32'hbf212ffa;
    11'd1827: sine = 32'hbf209394;
    11'd1828: sine = 32'hbf1ff6cc;
    11'd1829: sine = 32'hbf1f59a1;
    11'd1830: sine = 32'hbf1ebc13;
    11'd1831: sine = 32'hbf1e1e24;
    11'd1832: sine = 32'hbf1d7fd3;
    11'd1833: sine = 32'hbf1ce120;
    11'd1834: sine = 32'hbf1c420d;
    11'd1835: sine = 32'hbf1ba29a;
    11'd1836: sine = 32'hbf1b02c7;
    11'd1837: sine = 32'hbf1a6294;
    11'd1838: sine = 32'hbf19c202;
    11'd1839: sine = 32'hbf192111;
    11'd1840: sine = 32'hbf187fc1;
    11'd1841: sine = 32'hbf17de14;
    11'd1842: sine = 32'hbf173c08;
    11'd1843: sine = 32'hbf1699a0;
    11'd1844: sine = 32'hbf15f6da;
    11'd1845: sine = 32'hbf1553b9;
    11'd1846: sine = 32'hbf14b03b;
    11'd1847: sine = 32'hbf140c61;
    11'd1848: sine = 32'hbf13682c;
    11'd1849: sine = 32'hbf12c39c;
    11'd1850: sine = 32'hbf121eb1;
    11'd1851: sine = 32'hbf11796d;
    11'd1852: sine = 32'hbf10d3ce;
    11'd1853: sine = 32'hbf102dd6;
    11'd1854: sine = 32'hbf0f8786;
    11'd1855: sine = 32'hbf0ee0dd;
    11'd1856: sine = 32'hbf0e39db;
    11'd1857: sine = 32'hbf0d9282;
    11'd1858: sine = 32'hbf0cead2;
    11'd1859: sine = 32'hbf0c42ca;
    11'd1860: sine = 32'hbf0b9a6c;
    11'd1861: sine = 32'hbf0af1b9;
    11'd1862: sine = 32'hbf0a48af;
    11'd1863: sine = 32'hbf099f50;
    11'd1864: sine = 32'hbf08f59c;
    11'd1865: sine = 32'hbf084b94;
    11'd1866: sine = 32'hbf07a137;
    11'd1867: sine = 32'hbf06f687;
    11'd1868: sine = 32'hbf064b84;
    11'd1869: sine = 32'hbf05a02e;
    11'd1870: sine = 32'hbf04f485;
    11'd1871: sine = 32'hbf04488a;
    11'd1872: sine = 32'hbf039c3e;
    11'd1873: sine = 32'hbf02efa1;
    11'd1874: sine = 32'hbf0242b3;
    11'd1875: sine = 32'hbf019574;
    11'd1876: sine = 32'hbf00e7e6;
    11'd1877: sine = 32'hbf003a08;
    11'd1878: sine = 32'hbeff17b5;
    11'd1879: sine = 32'hbefdbabe;
    11'd1880: sine = 32'hbefc5d2a;
    11'd1881: sine = 32'hbefafefa;
    11'd1882: sine = 32'hbef9a030;
    11'd1883: sine = 32'hbef840cb;
    11'd1884: sine = 32'hbef6e0cd;
    11'd1885: sine = 32'hbef58038;
    11'd1886: sine = 32'hbef41f0a;
    11'd1887: sine = 32'hbef2bd46;
    11'd1888: sine = 32'hbef15aed;
    11'd1889: sine = 32'hbeeff7fe;
    11'd1890: sine = 32'hbeee947c;
    11'd1891: sine = 32'hbeed3066;
    11'd1892: sine = 32'hbeebcbbe;
    11'd1893: sine = 32'hbeea6684;
    11'd1894: sine = 32'hbee900ba;
    11'd1895: sine = 32'hbee79a60;
    11'd1896: sine = 32'hbee63378;
    11'd1897: sine = 32'hbee4cc01;
    11'd1898: sine = 32'hbee363fd;
    11'd1899: sine = 32'hbee1fb6d;
    11'd1900: sine = 32'hbee09252;
    11'd1901: sine = 32'hbedf28ac;
    11'd1902: sine = 32'hbeddbe7c;
    11'd1903: sine = 32'hbedc53c4;
    11'd1904: sine = 32'hbedae883;
    11'd1905: sine = 32'hbed97cbc;
    11'd1906: sine = 32'hbed8106e;
    11'd1907: sine = 32'hbed6a39c;
    11'd1908: sine = 32'hbed53644;
    11'd1909: sine = 32'hbed3c86a;
    11'd1910: sine = 32'hbed25a0c;
    11'd1911: sine = 32'hbed0eb2d;
    11'd1912: sine = 32'hbecf7bcd;
    11'd1913: sine = 32'hbece0bed;
    11'd1914: sine = 32'hbecc9b8e;
    11'd1915: sine = 32'hbecb2ab1;
    11'd1916: sine = 32'hbec9b956;
    11'd1917: sine = 32'hbec8477f;
    11'd1918: sine = 32'hbec6d52d;
    11'd1919: sine = 32'hbec5625f;
    11'd1920: sine = 32'hbec3ef18;
    11'd1921: sine = 32'hbec27b58;
    11'd1922: sine = 32'hbec10721;
    11'd1923: sine = 32'hbebf9272;
    11'd1924: sine = 32'hbebe1d4d;
    11'd1925: sine = 32'hbebca7b2;
    11'd1926: sine = 32'hbebb31a4;
    11'd1927: sine = 32'hbeb9bb21;
    11'd1928: sine = 32'hbeb8442d;
    11'd1929: sine = 32'hbeb6ccc6;
    11'd1930: sine = 32'hbeb554ef;
    11'd1931: sine = 32'hbeb3dca8;
    11'd1932: sine = 32'hbeb263f2;
    11'd1933: sine = 32'hbeb0eace;
    11'd1934: sine = 32'hbeaf713d;
    11'd1935: sine = 32'hbeadf740;
    11'd1936: sine = 32'hbeac7cd7;
    11'd1937: sine = 32'hbeab0204;
    11'd1938: sine = 32'hbea986c7;
    11'd1939: sine = 32'hbea80b22;
    11'd1940: sine = 32'hbea68f15;
    11'd1941: sine = 32'hbea512a2;
    11'd1942: sine = 32'hbea395c8;
    11'd1943: sine = 32'hbea2188a;
    11'd1944: sine = 32'hbea09ae8;
    11'd1945: sine = 32'hbe9f1ce3;
    11'd1946: sine = 32'hbe9d9e7b;
    11'd1947: sine = 32'hbe9c1fb2;
    11'd1948: sine = 32'hbe9aa089;
    11'd1949: sine = 32'hbe992101;
    11'd1950: sine = 32'hbe97a11a;
    11'd1951: sine = 32'hbe9620d6;
    11'd1952: sine = 32'hbe94a035;
    11'd1953: sine = 32'hbe931f38;
    11'd1954: sine = 32'hbe919de1;
    11'd1955: sine = 32'hbe901c2f;
    11'd1956: sine = 32'hbe8e9a25;
    11'd1957: sine = 32'hbe8d17c3;
    11'd1958: sine = 32'hbe8b950a;
    11'd1959: sine = 32'hbe8a11fb;
    11'd1960: sine = 32'hbe888e96;
    11'd1961: sine = 32'hbe870ade;
    11'd1962: sine = 32'hbe8586d2;
    11'd1963: sine = 32'hbe840274;
    11'd1964: sine = 32'hbe827dc4;
    11'd1965: sine = 32'hbe80f8c4;
    11'd1966: sine = 32'hbe7ee6e8;
    11'd1967: sine = 32'hbe7bdbab;
    11'd1968: sine = 32'hbe78cfd3;
    11'd1969: sine = 32'hbe75c361;
    11'd1970: sine = 32'hbe72b658;
    11'd1971: sine = 32'hbe6fa8b9;
    11'd1972: sine = 32'hbe6c9a86;
    11'd1973: sine = 32'hbe698bc1;
    11'd1974: sine = 32'hbe667c6c;
    11'd1975: sine = 32'hbe636c89;
    11'd1976: sine = 32'hbe605c1a;
    11'd1977: sine = 32'hbe5d4b20;
    11'd1978: sine = 32'hbe5a399e;
    11'd1979: sine = 32'hbe572795;
    11'd1980: sine = 32'hbe541508;
    11'd1981: sine = 32'hbe5101f8;
    11'd1982: sine = 32'hbe4dee66;
    11'd1983: sine = 32'hbe4ada56;
    11'd1984: sine = 32'hbe47c5c9;
    11'd1985: sine = 32'hbe44b0c0;
    11'd1986: sine = 32'hbe419b3e;
    11'd1987: sine = 32'hbe3e8545;
    11'd1988: sine = 32'hbe3b6ed6;
    11'd1989: sine = 32'hbe3857f3;
    11'd1990: sine = 32'hbe35409f;
    11'd1991: sine = 32'hbe3228db;
    11'd1992: sine = 32'hbe2f10a9;
    11'd1993: sine = 32'hbe2bf80b;
    11'd1994: sine = 32'hbe28df03;
    11'd1995: sine = 32'hbe25c593;
    11'd1996: sine = 32'hbe22abbc;
    11'd1997: sine = 32'hbe1f9182;
    11'd1998: sine = 32'hbe1c76e4;
    11'd1999: sine = 32'hbe195be7;
    11'd2000: sine = 32'hbe16408a;
    11'd2001: sine = 32'hbe1324d1;
    11'd2002: sine = 32'hbe1008be;
    11'd2003: sine = 32'hbe0cec51;
    11'd2004: sine = 32'hbe09cf8d;
    11'd2005: sine = 32'hbe06b275;
    11'd2006: sine = 32'hbe039509;
    11'd2007: sine = 32'hbe00774c;
    11'd2008: sine = 32'hbdfab281;
    11'd2009: sine = 32'hbdf475ce;
    11'd2010: sine = 32'hbdee3884;
    11'd2011: sine = 32'hbde7faa8;
    11'd2012: sine = 32'hbde1bc3c;
    11'd2013: sine = 32'hbddb7d45;
    11'd2014: sine = 32'hbdd53dc7;
    11'd2015: sine = 32'hbdcefdc5;
    11'd2016: sine = 32'hbdc8bd44;
    11'd2017: sine = 32'hbdc27c47;
    11'd2018: sine = 32'hbdbc3ad1;
    11'd2019: sine = 32'hbdb5f8e8;
    11'd2020: sine = 32'hbdafb68e;
    11'd2021: sine = 32'hbda973c8;
    11'd2022: sine = 32'hbda3309a;
    11'd2023: sine = 32'hbd9ced07;
    11'd2024: sine = 32'hbd96a913;
    11'd2025: sine = 32'hbd9064c2;
    11'd2026: sine = 32'hbd8a2018;
    11'd2027: sine = 32'hbd83db19;
    11'd2028: sine = 32'hbd7b2b90;
    11'd2029: sine = 32'hbd6ea054;
    11'd2030: sine = 32'hbd621485;
    11'd2031: sine = 32'hbd55882a;
    11'd2032: sine = 32'hbd48fb4c;
    11'd2033: sine = 32'hbd3c6df2;
    11'd2034: sine = 32'hbd2fe023;
    11'd2035: sine = 32'hbd2351e8;
    11'd2036: sine = 32'hbd16c348;
    11'd2037: sine = 32'hbd0a344b;
    11'd2038: sine = 32'hbcfb49f3;
    11'd2039: sine = 32'hbce22ab4;
    11'd2040: sine = 32'hbcc90ae9;
    11'd2041: sine = 32'hbcafeaa2;
    11'd2042: sine = 32'hbc96c9ef;
    11'd2043: sine = 32'hbc7b51be;
    11'd2044: sine = 32'hbc490f03;
    11'd2045: sine = 32'hbc16cbcb;
    11'd2046: sine = 32'hbbc9106e;
    11'd2047: sine = 32'hbb491192;
  endcase
end
endmodule
