`timescale 1ns/1ns
module sim_bldc
(input [2:0] hi,
 input [2:0] lo,
 output [15:0] current);



endmodule

