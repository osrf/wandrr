`timescale 1ns/1ns
module sine_table_11bit
(input c,
 input      [10:0] angle,
 output reg [31:0] sine);

always @(posedge c) begin
  case (angle)
    11'd0: sine = 32'h0;
    11'd1: sine = 32'h3e9d1452;
    11'd2: sine = 32'h3f1d1422;
    11'd3: sine = 32'h3f6b9dba;
    11'd4: sine = 32'h3f9d1360;
    11'd5: sine = 32'h3fc45783;
    11'd6: sine = 32'h3feb9b2c;
    11'd7: sine = 32'h40096f22;
    11'd8: sine = 32'h401d1059;
    11'd9: sine = 32'h4030b12f;
    11'd10: sine = 32'h40445199;
    11'd11: sine = 32'h4057f189;
    11'd12: sine = 32'h406b90f4;
    11'd13: sine = 32'h407f2fce;
    11'd14: sine = 32'h40896705;
    11'd15: sine = 32'h409335ce;
    11'd16: sine = 32'h409d043d;
    11'd17: sine = 32'h40a6d24b;
    11'd18: sine = 32'h40b09ff2;
    11'd19: sine = 32'h40ba6d2b;
    11'd20: sine = 32'h40c439f2;
    11'd21: sine = 32'h40ce0640;
    11'd22: sine = 32'h40d7d20f;
    11'd23: sine = 32'h40e19d58;
    11'd24: sine = 32'h40eb6817;
    11'd25: sine = 32'h40f53244;
    11'd26: sine = 32'h40fefbda;
    11'd27: sine = 32'h41046269;
    11'd28: sine = 32'h41094694;
    11'd29: sine = 32'h410e2a6a;
    11'd30: sine = 32'h41130de8;
    11'd31: sine = 32'h4117f10c;
    11'd32: sine = 32'h411cd3d2;
    11'd33: sine = 32'h4121b637;
    11'd34: sine = 32'h41269838;
    11'd35: sine = 32'h412b79d3;
    11'd36: sine = 32'h41305b04;
    11'd37: sine = 32'h41353bc8;
    11'd38: sine = 32'h413a1c1c;
    11'd39: sine = 32'h413efbfe;
    11'd40: sine = 32'h4143db69;
    11'd41: sine = 32'h4148ba5c;
    11'd42: sine = 32'h414d98d3;
    11'd43: sine = 32'h415276cb;
    11'd44: sine = 32'h41575442;
    11'd45: sine = 32'h415c3133;
    11'd46: sine = 32'h41610d9d;
    11'd47: sine = 32'h4165e97c;
    11'd48: sine = 32'h416ac4cd;
    11'd49: sine = 32'h416f9f8d;
    11'd50: sine = 32'h417479ba;
    11'd51: sine = 32'h41795350;
    11'd52: sine = 32'h417e2c4b;
    11'd53: sine = 32'h41818255;
    11'd54: sine = 32'h4183ee35;
    11'd55: sine = 32'h418659c3;
    11'd56: sine = 32'h4188c4ff;
    11'd57: sine = 32'h418b2fe6;
    11'd58: sine = 32'h418d9a77;
    11'd59: sine = 32'h419004b1;
    11'd60: sine = 32'h41926e92;
    11'd61: sine = 32'h4194d818;
    11'd62: sine = 32'h41974143;
    11'd63: sine = 32'h4199aa11;
    11'd64: sine = 32'h419c127f;
    11'd65: sine = 32'h419e7a8e;
    11'd66: sine = 32'h41a0e23b;
    11'd67: sine = 32'h41a34984;
    11'd68: sine = 32'h41a5b069;
    11'd69: sine = 32'h41a816e7;
    11'd70: sine = 32'h41aa7cfe;
    11'd71: sine = 32'h41ace2ac;
    11'd72: sine = 32'h41af47ef;
    11'd73: sine = 32'h41b1acc6;
    11'd74: sine = 32'h41b4112f;
    11'd75: sine = 32'h41b67529;
    11'd76: sine = 32'h41b8d8b3;
    11'd77: sine = 32'h41bb3bcb;
    11'd78: sine = 32'h41bd9e6f;
    11'd79: sine = 32'h41c0009e;
    11'd80: sine = 32'h41c26257;
    11'd81: sine = 32'h41c4c398;
    11'd82: sine = 32'h41c7245f;
    11'd83: sine = 32'h41c984ac;
    11'd84: sine = 32'h41cbe47c;
    11'd85: sine = 32'h41ce43cf;
    11'd86: sine = 32'h41d0a2a2;
    11'd87: sine = 32'h41d300f5;
    11'd88: sine = 32'h41d55ec6;
    11'd89: sine = 32'h41d7bc12;
    11'd90: sine = 32'h41da18da;
    11'd91: sine = 32'h41dc751c;
    11'd92: sine = 32'h41ded0d5;
    11'd93: sine = 32'h41e12c05;
    11'd94: sine = 32'h41e386aa;
    11'd95: sine = 32'h41e5e0c2;
    11'd96: sine = 32'h41e83a4d;
    11'd97: sine = 32'h41ea9349;
    11'd98: sine = 32'h41ecebb3;
    11'd99: sine = 32'h41ef438c;
    11'd100: sine = 32'h41f19ad1;
    11'd101: sine = 32'h41f3f181;
    11'd102: sine = 32'h41f6479b;
    11'd103: sine = 32'h41f89d1d;
    11'd104: sine = 32'h41faf205;
    11'd105: sine = 32'h41fd4652;
    11'd106: sine = 32'h41ff9a04;
    11'd107: sine = 32'h4200f68c;
    11'd108: sine = 32'h42021fc6;
    11'd109: sine = 32'h420348b0;
    11'd110: sine = 32'h42047149;
    11'd111: sine = 32'h42059990;
    11'd112: sine = 32'h4206c185;
    11'd113: sine = 32'h4207e927;
    11'd114: sine = 32'h42091075;
    11'd115: sine = 32'h420a376e;
    11'd116: sine = 32'h420b5e13;
    11'd117: sine = 32'h420c8461;
    11'd118: sine = 32'h420daa58;
    11'd119: sine = 32'h420ecff8;
    11'd120: sine = 32'h420ff540;
    11'd121: sine = 32'h42111a30;
    11'd122: sine = 32'h42123ec5;
    11'd123: sine = 32'h42136301;
    11'd124: sine = 32'h421486e1;
    11'd125: sine = 32'h4215aa66;
    11'd126: sine = 32'h4216cd8f;
    11'd127: sine = 32'h4217f05b;
    11'd128: sine = 32'h421912c8;
    11'd129: sine = 32'h421a34d8;
    11'd130: sine = 32'h421b5688;
    11'd131: sine = 32'h421c77d9;
    11'd132: sine = 32'h421d98c9;
    11'd133: sine = 32'h421eb958;
    11'd134: sine = 32'h421fd984;
    11'd135: sine = 32'h4220f94f;
    11'd136: sine = 32'h422218b6;
    11'd137: sine = 32'h422337b9;
    11'd138: sine = 32'h42245657;
    11'd139: sine = 32'h42257490;
    11'd140: sine = 32'h42269263;
    11'd141: sine = 32'h4227afcf;
    11'd142: sine = 32'h4228ccd4;
    11'd143: sine = 32'h4229e970;
    11'd144: sine = 32'h422b05a4;
    11'd145: sine = 32'h422c216e;
    11'd146: sine = 32'h422d3cce;
    11'd147: sine = 32'h422e57c4;
    11'd148: sine = 32'h422f724d;
    11'd149: sine = 32'h42308c6b;
    11'd150: sine = 32'h4231a61b;
    11'd151: sine = 32'h4232bf5e;
    11'd152: sine = 32'h4233d833;
    11'd153: sine = 32'h4234f099;
    11'd154: sine = 32'h4236088f;
    11'd155: sine = 32'h42372015;
    11'd156: sine = 32'h4238372a;
    11'd157: sine = 32'h42394dcd;
    11'd158: sine = 32'h423a63fe;
    11'd159: sine = 32'h423b79bc;
    11'd160: sine = 32'h423c8f06;
    11'd161: sine = 32'h423da3dc;
    11'd162: sine = 32'h423eb83e;
    11'd163: sine = 32'h423fcc29;
    11'd164: sine = 32'h4240df9e;
    11'd165: sine = 32'h4241f29c;
    11'd166: sine = 32'h42430523;
    11'd167: sine = 32'h42441731;
    11'd168: sine = 32'h424528c6;
    11'd169: sine = 32'h424639e2;
    11'd170: sine = 32'h42474a83;
    11'd171: sine = 32'h42485aaa;
    11'd172: sine = 32'h42496a54;
    11'd173: sine = 32'h424a7983;
    11'd174: sine = 32'h424b8835;
    11'd175: sine = 32'h424c9669;
    11'd176: sine = 32'h424da41f;
    11'd177: sine = 32'h424eb156;
    11'd178: sine = 32'h424fbe0d;
    11'd179: sine = 32'h4250ca45;
    11'd180: sine = 32'h4251d5fc;
    11'd181: sine = 32'h4252e131;
    11'd182: sine = 32'h4253ebe4;
    11'd183: sine = 32'h4254f614;
    11'd184: sine = 32'h4255ffc1;
    11'd185: sine = 32'h425708ea;
    11'd186: sine = 32'h4258118f;
    11'd187: sine = 32'h425919ae;
    11'd188: sine = 32'h425a2147;
    11'd189: sine = 32'h425b285a;
    11'd190: sine = 32'h425c2ee5;
    11'd191: sine = 32'h425d34e9;
    11'd192: sine = 32'h425e3a64;
    11'd193: sine = 32'h425f3f56;
    11'd194: sine = 32'h426043bf;
    11'd195: sine = 32'h4261479d;
    11'd196: sine = 32'h42624af0;
    11'd197: sine = 32'h42634db7;
    11'd198: sine = 32'h42644ff3;
    11'd199: sine = 32'h426551a1;
    11'd200: sine = 32'h426652c2;
    11'd201: sine = 32'h42675355;
    11'd202: sine = 32'h42685359;
    11'd203: sine = 32'h426952ce;
    11'd204: sine = 32'h426a51b3;
    11'd205: sine = 32'h426b5008;
    11'd206: sine = 32'h426c4dcb;
    11'd207: sine = 32'h426d4afc;
    11'd208: sine = 32'h426e479c;
    11'd209: sine = 32'h426f43a8;
    11'd210: sine = 32'h42703f20;
    11'd211: sine = 32'h42713a05;
    11'd212: sine = 32'h42723454;
    11'd213: sine = 32'h42732e0f;
    11'd214: sine = 32'h42742733;
    11'd215: sine = 32'h42751fc0;
    11'd216: sine = 32'h427617b7;
    11'd217: sine = 32'h42770f15;
    11'd218: sine = 32'h427805dc;
    11'd219: sine = 32'h4278fc09;
    11'd220: sine = 32'h4279f19c;
    11'd221: sine = 32'h427ae696;
    11'd222: sine = 32'h427bdaf4;
    11'd223: sine = 32'h427cceb8;
    11'd224: sine = 32'h427dc1df;
    11'd225: sine = 32'h427eb46a;
    11'd226: sine = 32'h427fa658;
    11'd227: sine = 32'h42804bd4;
    11'd228: sine = 32'h4280c42d;
    11'd229: sine = 32'h42813c36;
    11'd230: sine = 32'h4281b3f0;
    11'd231: sine = 32'h42822b5a;
    11'd232: sine = 32'h4282a273;
    11'd233: sine = 32'h4283193c;
    11'd234: sine = 32'h42838fb4;
    11'd235: sine = 32'h428405db;
    11'd236: sine = 32'h42847bb0;
    11'd237: sine = 32'h4284f134;
    11'd238: sine = 32'h42856665;
    11'd239: sine = 32'h4285db45;
    11'd240: sine = 32'h42864fd1;
    11'd241: sine = 32'h4286c40b;
    11'd242: sine = 32'h428737f2;
    11'd243: sine = 32'h4287ab86;
    11'd244: sine = 32'h42881ec5;
    11'd245: sine = 32'h428891b1;
    11'd246: sine = 32'h42890449;
    11'd247: sine = 32'h4289768c;
    11'd248: sine = 32'h4289e87a;
    11'd249: sine = 32'h428a5a13;
    11'd250: sine = 32'h428acb57;
    11'd251: sine = 32'h428b3c45;
    11'd252: sine = 32'h428bacdd;
    11'd253: sine = 32'h428c1d1f;
    11'd254: sine = 32'h428c8d0b;
    11'd255: sine = 32'h428cfca0;
    11'd256: sine = 32'h428d6bde;
    11'd257: sine = 32'h428ddac5;
    11'd258: sine = 32'h428e4954;
    11'd259: sine = 32'h428eb78b;
    11'd260: sine = 32'h428f256b;
    11'd261: sine = 32'h428f92f2;
    11'd262: sine = 32'h42900021;
    11'd263: sine = 32'h42906cf7;
    11'd264: sine = 32'h4290d973;
    11'd265: sine = 32'h42914597;
    11'd266: sine = 32'h4291b160;
    11'd267: sine = 32'h42921cd0;
    11'd268: sine = 32'h429287e6;
    11'd269: sine = 32'h4292f2a1;
    11'd270: sine = 32'h42935d02;
    11'd271: sine = 32'h4293c708;
    11'd272: sine = 32'h429430b2;
    11'd273: sine = 32'h42949a02;
    11'd274: sine = 32'h429502f5;
    11'd275: sine = 32'h42956b8d;
    11'd276: sine = 32'h4295d3c8;
    11'd277: sine = 32'h42963ba7;
    11'd278: sine = 32'h4296a32a;
    11'd279: sine = 32'h42970a4f;
    11'd280: sine = 32'h42977118;
    11'd281: sine = 32'h4297d783;
    11'd282: sine = 32'h42983d90;
    11'd283: sine = 32'h4298a33f;
    11'd284: sine = 32'h42990890;
    11'd285: sine = 32'h42996d83;
    11'd286: sine = 32'h4299d217;
    11'd287: sine = 32'h429a364c;
    11'd288: sine = 32'h429a9a22;
    11'd289: sine = 32'h429afd99;
    11'd290: sine = 32'h429b60b0;
    11'd291: sine = 32'h429bc368;
    11'd292: sine = 32'h429c25bf;
    11'd293: sine = 32'h429c87b6;
    11'd294: sine = 32'h429ce94c;
    11'd295: sine = 32'h429d4a82;
    11'd296: sine = 32'h429dab56;
    11'd297: sine = 32'h429e0bc9;
    11'd298: sine = 32'h429e6bdb;
    11'd299: sine = 32'h429ecb8b;
    11'd300: sine = 32'h429f2ad9;
    11'd301: sine = 32'h429f89c5;
    11'd302: sine = 32'h429fe84f;
    11'd303: sine = 32'h42a04676;
    11'd304: sine = 32'h42a0a43a;
    11'd305: sine = 32'h42a1019b;
    11'd306: sine = 32'h42a15e98;
    11'd307: sine = 32'h42a1bb32;
    11'd308: sine = 32'h42a21768;
    11'd309: sine = 32'h42a2733b;
    11'd310: sine = 32'h42a2cea9;
    11'd311: sine = 32'h42a329b3;
    11'd312: sine = 32'h42a38458;
    11'd313: sine = 32'h42a3de98;
    11'd314: sine = 32'h42a43873;
    11'd315: sine = 32'h42a491e9;
    11'd316: sine = 32'h42a4eaf9;
    11'd317: sine = 32'h42a543a3;
    11'd318: sine = 32'h42a59be8;
    11'd319: sine = 32'h42a5f3c6;
    11'd320: sine = 32'h42a64b3e;
    11'd321: sine = 32'h42a6a250;
    11'd322: sine = 32'h42a6f8fb;
    11'd323: sine = 32'h42a74f3e;
    11'd324: sine = 32'h42a7a51b;
    11'd325: sine = 32'h42a7fa90;
    11'd326: sine = 32'h42a84f9d;
    11'd327: sine = 32'h42a8a443;
    11'd328: sine = 32'h42a8f881;
    11'd329: sine = 32'h42a94c56;
    11'd330: sine = 32'h42a99fc3;
    11'd331: sine = 32'h42a9f2c7;
    11'd332: sine = 32'h42aa4563;
    11'd333: sine = 32'h42aa9795;
    11'd334: sine = 32'h42aae95e;
    11'd335: sine = 32'h42ab3abe;
    11'd336: sine = 32'h42ab8bb4;
    11'd337: sine = 32'h42abdc41;
    11'd338: sine = 32'h42ac2c63;
    11'd339: sine = 32'h42ac7c1b;
    11'd340: sine = 32'h42accb69;
    11'd341: sine = 32'h42ad1a4c;
    11'd342: sine = 32'h42ad68c4;
    11'd343: sine = 32'h42adb6d2;
    11'd344: sine = 32'h42ae0474;
    11'd345: sine = 32'h42ae51ab;
    11'd346: sine = 32'h42ae9e76;
    11'd347: sine = 32'h42aeead6;
    11'd348: sine = 32'h42af36ca;
    11'd349: sine = 32'h42af8252;
    11'd350: sine = 32'h42afcd6d;
    11'd351: sine = 32'h42b0181c;
    11'd352: sine = 32'h42b0625e;
    11'd353: sine = 32'h42b0ac34;
    11'd354: sine = 32'h42b0f59c;
    11'd355: sine = 32'h42b13e98;
    11'd356: sine = 32'h42b18726;
    11'd357: sine = 32'h42b1cf46;
    11'd358: sine = 32'h42b216f9;
    11'd359: sine = 32'h42b25e3e;
    11'd360: sine = 32'h42b2a515;
    11'd361: sine = 32'h42b2eb7e;
    11'd362: sine = 32'h42b33179;
    11'd363: sine = 32'h42b37705;
    11'd364: sine = 32'h42b3bc22;
    11'd365: sine = 32'h42b400d0;
    11'd366: sine = 32'h42b4450f;
    11'd367: sine = 32'h42b488e0;
    11'd368: sine = 32'h42b4cc40;
    11'd369: sine = 32'h42b50f32;
    11'd370: sine = 32'h42b551b3;
    11'd371: sine = 32'h42b593c5;
    11'd372: sine = 32'h42b5d566;
    11'd373: sine = 32'h42b61698;
    11'd374: sine = 32'h42b65759;
    11'd375: sine = 32'h42b697aa;
    11'd376: sine = 32'h42b6d78a;
    11'd377: sine = 32'h42b716f9;
    11'd378: sine = 32'h42b755f8;
    11'd379: sine = 32'h42b79485;
    11'd380: sine = 32'h42b7d2a1;
    11'd381: sine = 32'h42b8104c;
    11'd382: sine = 32'h42b84d85;
    11'd383: sine = 32'h42b88a4c;
    11'd384: sine = 32'h42b8c6a2;
    11'd385: sine = 32'h42b90285;
    11'd386: sine = 32'h42b93df7;
    11'd387: sine = 32'h42b978f6;
    11'd388: sine = 32'h42b9b383;
    11'd389: sine = 32'h42b9ed9d;
    11'd390: sine = 32'h42ba2745;
    11'd391: sine = 32'h42ba6079;
    11'd392: sine = 32'h42ba993b;
    11'd393: sine = 32'h42bad18a;
    11'd394: sine = 32'h42bb0965;
    11'd395: sine = 32'h42bb40cd;
    11'd396: sine = 32'h42bb77c2;
    11'd397: sine = 32'h42bbae43;
    11'd398: sine = 32'h42bbe450;
    11'd399: sine = 32'h42bc19e9;
    11'd400: sine = 32'h42bc4f0e;
    11'd401: sine = 32'h42bc83bf;
    11'd402: sine = 32'h42bcb7fc;
    11'd403: sine = 32'h42bcebc4;
    11'd404: sine = 32'h42bd1f18;
    11'd405: sine = 32'h42bd51f7;
    11'd406: sine = 32'h42bd8462;
    11'd407: sine = 32'h42bdb657;
    11'd408: sine = 32'h42bde7d8;
    11'd409: sine = 32'h42be18e3;
    11'd410: sine = 32'h42be4979;
    11'd411: sine = 32'h42be799a;
    11'd412: sine = 32'h42bea945;
    11'd413: sine = 32'h42bed87a;
    11'd414: sine = 32'h42bf073a;
    11'd415: sine = 32'h42bf3584;
    11'd416: sine = 32'h42bf6358;
    11'd417: sine = 32'h42bf90b6;
    11'd418: sine = 32'h42bfbd9e;
    11'd419: sine = 32'h42bfea10;
    11'd420: sine = 32'h42c0160b;
    11'd421: sine = 32'h42c04190;
    11'd422: sine = 32'h42c06c9e;
    11'd423: sine = 32'h42c09735;
    11'd424: sine = 32'h42c0c156;
    11'd425: sine = 32'h42c0eaff;
    11'd426: sine = 32'h42c11432;
    11'd427: sine = 32'h42c13cee;
    11'd428: sine = 32'h42c16532;
    11'd429: sine = 32'h42c18cff;
    11'd430: sine = 32'h42c1b455;
    11'd431: sine = 32'h42c1db33;
    11'd432: sine = 32'h42c2019a;
    11'd433: sine = 32'h42c22789;
    11'd434: sine = 32'h42c24d00;
    11'd435: sine = 32'h42c271ff;
    11'd436: sine = 32'h42c29686;
    11'd437: sine = 32'h42c2ba96;
    11'd438: sine = 32'h42c2de2d;
    11'd439: sine = 32'h42c3014c;
    11'd440: sine = 32'h42c323f3;
    11'd441: sine = 32'h42c34621;
    11'd442: sine = 32'h42c367d7;
    11'd443: sine = 32'h42c38915;
    11'd444: sine = 32'h42c3a9d9;
    11'd445: sine = 32'h42c3ca25;
    11'd446: sine = 32'h42c3e9f9;
    11'd447: sine = 32'h42c40953;
    11'd448: sine = 32'h42c42835;
    11'd449: sine = 32'h42c4469d;
    11'd450: sine = 32'h42c4648d;
    11'd451: sine = 32'h42c48203;
    11'd452: sine = 32'h42c49f00;
    11'd453: sine = 32'h42c4bb84;
    11'd454: sine = 32'h42c4d78e;
    11'd455: sine = 32'h42c4f320;
    11'd456: sine = 32'h42c50e37;
    11'd457: sine = 32'h42c528d5;
    11'd458: sine = 32'h42c542f9;
    11'd459: sine = 32'h42c55ca4;
    11'd460: sine = 32'h42c575d5;
    11'd461: sine = 32'h42c58e8c;
    11'd462: sine = 32'h42c5a6ca;
    11'd463: sine = 32'h42c5be8d;
    11'd464: sine = 32'h42c5d5d6;
    11'd465: sine = 32'h42c5eca6;
    11'd466: sine = 32'h42c602fb;
    11'd467: sine = 32'h42c618d6;
    11'd468: sine = 32'h42c62e37;
    11'd469: sine = 32'h42c6431e;
    11'd470: sine = 32'h42c6578a;
    11'd471: sine = 32'h42c66b7c;
    11'd472: sine = 32'h42c67ef4;
    11'd473: sine = 32'h42c691f1;
    11'd474: sine = 32'h42c6a474;
    11'd475: sine = 32'h42c6b67c;
    11'd476: sine = 32'h42c6c809;
    11'd477: sine = 32'h42c6d91c;
    11'd478: sine = 32'h42c6e9b5;
    11'd479: sine = 32'h42c6f9d2;
    11'd480: sine = 32'h42c70975;
    11'd481: sine = 32'h42c7189d;
    11'd482: sine = 32'h42c7274b;
    11'd483: sine = 32'h42c7357d;
    11'd484: sine = 32'h42c74335;
    11'd485: sine = 32'h42c75071;
    11'd486: sine = 32'h42c75d33;
    11'd487: sine = 32'h42c7697a;
    11'd488: sine = 32'h42c77545;
    11'd489: sine = 32'h42c78096;
    11'd490: sine = 32'h42c78b6c;
    11'd491: sine = 32'h42c795c6;
    11'd492: sine = 32'h42c79fa6;
    11'd493: sine = 32'h42c7a90a;
    11'd494: sine = 32'h42c7b1f3;
    11'd495: sine = 32'h42c7ba61;
    11'd496: sine = 32'h42c7c254;
    11'd497: sine = 32'h42c7c9cb;
    11'd498: sine = 32'h42c7d0c8;
    11'd499: sine = 32'h42c7d749;
    11'd500: sine = 32'h42c7dd4e;
    11'd501: sine = 32'h42c7e2d9;
    11'd502: sine = 32'h42c7e7e8;
    11'd503: sine = 32'h42c7ec7c;
    11'd504: sine = 32'h42c7f094;
    11'd505: sine = 32'h42c7f432;
    11'd506: sine = 32'h42c7f753;
    11'd507: sine = 32'h42c7f9fa;
    11'd508: sine = 32'h42c7fc25;
    11'd509: sine = 32'h42c7fdd5;
    11'd510: sine = 32'h42c7ff09;
    11'd511: sine = 32'h42c7ffc2;
    11'd512: sine = 32'h42c80000;
    11'd513: sine = 32'h42c7ffc2;
    11'd514: sine = 32'h42c7ff09;
    11'd515: sine = 32'h42c7fdd5;
    11'd516: sine = 32'h42c7fc25;
    11'd517: sine = 32'h42c7f9fa;
    11'd518: sine = 32'h42c7f753;
    11'd519: sine = 32'h42c7f432;
    11'd520: sine = 32'h42c7f094;
    11'd521: sine = 32'h42c7ec7c;
    11'd522: sine = 32'h42c7e7e8;
    11'd523: sine = 32'h42c7e2d9;
    11'd524: sine = 32'h42c7dd4e;
    11'd525: sine = 32'h42c7d749;
    11'd526: sine = 32'h42c7d0c8;
    11'd527: sine = 32'h42c7c9cb;
    11'd528: sine = 32'h42c7c254;
    11'd529: sine = 32'h42c7ba61;
    11'd530: sine = 32'h42c7b1f3;
    11'd531: sine = 32'h42c7a90a;
    11'd532: sine = 32'h42c79fa6;
    11'd533: sine = 32'h42c795c6;
    11'd534: sine = 32'h42c78b6c;
    11'd535: sine = 32'h42c78096;
    11'd536: sine = 32'h42c77546;
    11'd537: sine = 32'h42c7697a;
    11'd538: sine = 32'h42c75d33;
    11'd539: sine = 32'h42c75071;
    11'd540: sine = 32'h42c74335;
    11'd541: sine = 32'h42c7357d;
    11'd542: sine = 32'h42c7274b;
    11'd543: sine = 32'h42c7189d;
    11'd544: sine = 32'h42c70975;
    11'd545: sine = 32'h42c6f9d2;
    11'd546: sine = 32'h42c6e9b5;
    11'd547: sine = 32'h42c6d91c;
    11'd548: sine = 32'h42c6c809;
    11'd549: sine = 32'h42c6b67c;
    11'd550: sine = 32'h42c6a474;
    11'd551: sine = 32'h42c691f1;
    11'd552: sine = 32'h42c67ef4;
    11'd553: sine = 32'h42c66b7c;
    11'd554: sine = 32'h42c6578a;
    11'd555: sine = 32'h42c6431e;
    11'd556: sine = 32'h42c62e37;
    11'd557: sine = 32'h42c618d6;
    11'd558: sine = 32'h42c602fb;
    11'd559: sine = 32'h42c5eca6;
    11'd560: sine = 32'h42c5d5d6;
    11'd561: sine = 32'h42c5be8d;
    11'd562: sine = 32'h42c5a6ca;
    11'd563: sine = 32'h42c58e8c;
    11'd564: sine = 32'h42c575d5;
    11'd565: sine = 32'h42c55ca4;
    11'd566: sine = 32'h42c542fa;
    11'd567: sine = 32'h42c528d5;
    11'd568: sine = 32'h42c50e37;
    11'd569: sine = 32'h42c4f320;
    11'd570: sine = 32'h42c4d78f;
    11'd571: sine = 32'h42c4bb84;
    11'd572: sine = 32'h42c49f00;
    11'd573: sine = 32'h42c48203;
    11'd574: sine = 32'h42c4648d;
    11'd575: sine = 32'h42c4469d;
    11'd576: sine = 32'h42c42835;
    11'd577: sine = 32'h42c40953;
    11'd578: sine = 32'h42c3e9f9;
    11'd579: sine = 32'h42c3ca26;
    11'd580: sine = 32'h42c3a9da;
    11'd581: sine = 32'h42c38915;
    11'd582: sine = 32'h42c367d7;
    11'd583: sine = 32'h42c34621;
    11'd584: sine = 32'h42c323f3;
    11'd585: sine = 32'h42c3014c;
    11'd586: sine = 32'h42c2de2d;
    11'd587: sine = 32'h42c2ba96;
    11'd588: sine = 32'h42c29687;
    11'd589: sine = 32'h42c271ff;
    11'd590: sine = 32'h42c24d00;
    11'd591: sine = 32'h42c22789;
    11'd592: sine = 32'h42c2019a;
    11'd593: sine = 32'h42c1db33;
    11'd594: sine = 32'h42c1b455;
    11'd595: sine = 32'h42c18cff;
    11'd596: sine = 32'h42c16532;
    11'd597: sine = 32'h42c13cee;
    11'd598: sine = 32'h42c11432;
    11'd599: sine = 32'h42c0eaff;
    11'd600: sine = 32'h42c0c156;
    11'd601: sine = 32'h42c09735;
    11'd602: sine = 32'h42c06c9e;
    11'd603: sine = 32'h42c04190;
    11'd604: sine = 32'h42c0160b;
    11'd605: sine = 32'h42bfea10;
    11'd606: sine = 32'h42bfbd9e;
    11'd607: sine = 32'h42bf90b6;
    11'd608: sine = 32'h42bf6358;
    11'd609: sine = 32'h42bf3584;
    11'd610: sine = 32'h42bf073a;
    11'd611: sine = 32'h42bed87b;
    11'd612: sine = 32'h42bea945;
    11'd613: sine = 32'h42be799a;
    11'd614: sine = 32'h42be4979;
    11'd615: sine = 32'h42be18e3;
    11'd616: sine = 32'h42bde7d8;
    11'd617: sine = 32'h42bdb657;
    11'd618: sine = 32'h42bd8462;
    11'd619: sine = 32'h42bd51f8;
    11'd620: sine = 32'h42bd1f18;
    11'd621: sine = 32'h42bcebc5;
    11'd622: sine = 32'h42bcb7fc;
    11'd623: sine = 32'h42bc83c0;
    11'd624: sine = 32'h42bc4f0f;
    11'd625: sine = 32'h42bc19e9;
    11'd626: sine = 32'h42bbe450;
    11'd627: sine = 32'h42bbae43;
    11'd628: sine = 32'h42bb77c2;
    11'd629: sine = 32'h42bb40ce;
    11'd630: sine = 32'h42bb0965;
    11'd631: sine = 32'h42bad18a;
    11'd632: sine = 32'h42ba993b;
    11'd633: sine = 32'h42ba607a;
    11'd634: sine = 32'h42ba2745;
    11'd635: sine = 32'h42b9ed9d;
    11'd636: sine = 32'h42b9b383;
    11'd637: sine = 32'h42b978f6;
    11'd638: sine = 32'h42b93df7;
    11'd639: sine = 32'h42b90286;
    11'd640: sine = 32'h42b8c6a2;
    11'd641: sine = 32'h42b88a4c;
    11'd642: sine = 32'h42b84d85;
    11'd643: sine = 32'h42b8104c;
    11'd644: sine = 32'h42b7d2a1;
    11'd645: sine = 32'h42b79485;
    11'd646: sine = 32'h42b755f8;
    11'd647: sine = 32'h42b716fa;
    11'd648: sine = 32'h42b6d78a;
    11'd649: sine = 32'h42b697aa;
    11'd650: sine = 32'h42b65759;
    11'd651: sine = 32'h42b61698;
    11'd652: sine = 32'h42b5d567;
    11'd653: sine = 32'h42b593c5;
    11'd654: sine = 32'h42b551b3;
    11'd655: sine = 32'h42b50f32;
    11'd656: sine = 32'h42b4cc41;
    11'd657: sine = 32'h42b488e0;
    11'd658: sine = 32'h42b44510;
    11'd659: sine = 32'h42b400d0;
    11'd660: sine = 32'h42b3bc22;
    11'd661: sine = 32'h42b37705;
    11'd662: sine = 32'h42b33179;
    11'd663: sine = 32'h42b2eb7f;
    11'd664: sine = 32'h42b2a516;
    11'd665: sine = 32'h42b25e3f;
    11'd666: sine = 32'h42b216fa;
    11'd667: sine = 32'h42b1cf47;
    11'd668: sine = 32'h42b18726;
    11'd669: sine = 32'h42b13e98;
    11'd670: sine = 32'h42b0f59d;
    11'd671: sine = 32'h42b0ac34;
    11'd672: sine = 32'h42b0625f;
    11'd673: sine = 32'h42b0181c;
    11'd674: sine = 32'h42afcd6d;
    11'd675: sine = 32'h42af8252;
    11'd676: sine = 32'h42af36ca;
    11'd677: sine = 32'h42aeead6;
    11'd678: sine = 32'h42ae9e77;
    11'd679: sine = 32'h42ae51ab;
    11'd680: sine = 32'h42ae0474;
    11'd681: sine = 32'h42adb6d2;
    11'd682: sine = 32'h42ad68c5;
    11'd683: sine = 32'h42ad1a4c;
    11'd684: sine = 32'h42accb69;
    11'd685: sine = 32'h42ac7c1c;
    11'd686: sine = 32'h42ac2c63;
    11'd687: sine = 32'h42abdc41;
    11'd688: sine = 32'h42ab8bb5;
    11'd689: sine = 32'h42ab3abf;
    11'd690: sine = 32'h42aae95f;
    11'd691: sine = 32'h42aa9795;
    11'd692: sine = 32'h42aa4563;
    11'd693: sine = 32'h42a9f2c8;
    11'd694: sine = 32'h42a99fc3;
    11'd695: sine = 32'h42a94c56;
    11'd696: sine = 32'h42a8f881;
    11'd697: sine = 32'h42a8a443;
    11'd698: sine = 32'h42a84f9e;
    11'd699: sine = 32'h42a7fa90;
    11'd700: sine = 32'h42a7a51b;
    11'd701: sine = 32'h42a74f3f;
    11'd702: sine = 32'h42a6f8fb;
    11'd703: sine = 32'h42a6a250;
    11'd704: sine = 32'h42a64b3f;
    11'd705: sine = 32'h42a5f3c7;
    11'd706: sine = 32'h42a59be8;
    11'd707: sine = 32'h42a543a4;
    11'd708: sine = 32'h42a4eaf9;
    11'd709: sine = 32'h42a491e9;
    11'd710: sine = 32'h42a43873;
    11'd711: sine = 32'h42a3de98;
    11'd712: sine = 32'h42a38458;
    11'd713: sine = 32'h42a329b3;
    11'd714: sine = 32'h42a2cea9;
    11'd715: sine = 32'h42a2733b;
    11'd716: sine = 32'h42a21769;
    11'd717: sine = 32'h42a1bb33;
    11'd718: sine = 32'h42a15e99;
    11'd719: sine = 32'h42a1019b;
    11'd720: sine = 32'h42a0a43a;
    11'd721: sine = 32'h42a04676;
    11'd722: sine = 32'h429fe84f;
    11'd723: sine = 32'h429f89c6;
    11'd724: sine = 32'h429f2ada;
    11'd725: sine = 32'h429ecb8c;
    11'd726: sine = 32'h429e6bdc;
    11'd727: sine = 32'h429e0bca;
    11'd728: sine = 32'h429dab57;
    11'd729: sine = 32'h429d4a82;
    11'd730: sine = 32'h429ce94d;
    11'd731: sine = 32'h429c87b6;
    11'd732: sine = 32'h429c25bf;
    11'd733: sine = 32'h429bc368;
    11'd734: sine = 32'h429b60b1;
    11'd735: sine = 32'h429afd9a;
    11'd736: sine = 32'h429a9a23;
    11'd737: sine = 32'h429a364d;
    11'd738: sine = 32'h4299d218;
    11'd739: sine = 32'h42996d83;
    11'd740: sine = 32'h42990891;
    11'd741: sine = 32'h4298a340;
    11'd742: sine = 32'h42983d90;
    11'd743: sine = 32'h4297d783;
    11'd744: sine = 32'h42977118;
    11'd745: sine = 32'h42970a50;
    11'd746: sine = 32'h4296a32a;
    11'd747: sine = 32'h42963ba8;
    11'd748: sine = 32'h4295d3c9;
    11'd749: sine = 32'h42956b8d;
    11'd750: sine = 32'h429502f6;
    11'd751: sine = 32'h42949a02;
    11'd752: sine = 32'h429430b3;
    11'd753: sine = 32'h4293c708;
    11'd754: sine = 32'h42935d02;
    11'd755: sine = 32'h4292f2a2;
    11'd756: sine = 32'h429287e6;
    11'd757: sine = 32'h42921cd1;
    11'd758: sine = 32'h4291b161;
    11'd759: sine = 32'h42914597;
    11'd760: sine = 32'h4290d974;
    11'd761: sine = 32'h42906cf7;
    11'd762: sine = 32'h42900021;
    11'd763: sine = 32'h428f92f3;
    11'd764: sine = 32'h428f256b;
    11'd765: sine = 32'h428eb78c;
    11'd766: sine = 32'h428e4954;
    11'd767: sine = 32'h428ddac5;
    11'd768: sine = 32'h428d6bde;
    11'd769: sine = 32'h428cfca0;
    11'd770: sine = 32'h428c8d0b;
    11'd771: sine = 32'h428c1d20;
    11'd772: sine = 32'h428bacde;
    11'd773: sine = 32'h428b3c45;
    11'd774: sine = 32'h428acb57;
    11'd775: sine = 32'h428a5a13;
    11'd776: sine = 32'h4289e87a;
    11'd777: sine = 32'h4289768c;
    11'd778: sine = 32'h42890449;
    11'd779: sine = 32'h428891b2;
    11'd780: sine = 32'h42881ec6;
    11'd781: sine = 32'h4287ab86;
    11'd782: sine = 32'h428737f3;
    11'd783: sine = 32'h4286c40c;
    11'd784: sine = 32'h42864fd2;
    11'd785: sine = 32'h4285db45;
    11'd786: sine = 32'h42856666;
    11'd787: sine = 32'h4284f134;
    11'd788: sine = 32'h42847bb0;
    11'd789: sine = 32'h428405db;
    11'd790: sine = 32'h42838fb4;
    11'd791: sine = 32'h4283193c;
    11'd792: sine = 32'h4282a273;
    11'd793: sine = 32'h42822b5a;
    11'd794: sine = 32'h4281b3f0;
    11'd795: sine = 32'h42813c37;
    11'd796: sine = 32'h4280c42d;
    11'd797: sine = 32'h42804bd4;
    11'd798: sine = 32'h427fa659;
    11'd799: sine = 32'h427eb46b;
    11'd800: sine = 32'h427dc1e0;
    11'd801: sine = 32'h427cceb9;
    11'd802: sine = 32'h427bdaf6;
    11'd803: sine = 32'h427ae697;
    11'd804: sine = 32'h4279f19d;
    11'd805: sine = 32'h4278fc0a;
    11'd806: sine = 32'h427805dd;
    11'd807: sine = 32'h42770f16;
    11'd808: sine = 32'h427617b8;
    11'd809: sine = 32'h42751fc2;
    11'd810: sine = 32'h42742734;
    11'd811: sine = 32'h42732e10;
    11'd812: sine = 32'h42723456;
    11'd813: sine = 32'h42713a06;
    11'd814: sine = 32'h42703f22;
    11'd815: sine = 32'h426f43a9;
    11'd816: sine = 32'h426e479d;
    11'd817: sine = 32'h426d4afe;
    11'd818: sine = 32'h426c4dcc;
    11'd819: sine = 32'h426b5009;
    11'd820: sine = 32'h426a51b4;
    11'd821: sine = 32'h426952cf;
    11'd822: sine = 32'h4268535a;
    11'd823: sine = 32'h42675356;
    11'd824: sine = 32'h426652c3;
    11'd825: sine = 32'h426551a2;
    11'd826: sine = 32'h42644ff4;
    11'd827: sine = 32'h42634db8;
    11'd828: sine = 32'h42624af1;
    11'd829: sine = 32'h4261479e;
    11'd830: sine = 32'h426043c0;
    11'd831: sine = 32'h425f3f57;
    11'd832: sine = 32'h425e3a65;
    11'd833: sine = 32'h425d34ea;
    11'd834: sine = 32'h425c2ee6;
    11'd835: sine = 32'h425b285b;
    11'd836: sine = 32'h425a2148;
    11'd837: sine = 32'h425919af;
    11'd838: sine = 32'h42581190;
    11'd839: sine = 32'h425708ec;
    11'd840: sine = 32'h4255ffc3;
    11'd841: sine = 32'h4254f616;
    11'd842: sine = 32'h4253ebe5;
    11'd843: sine = 32'h4252e132;
    11'd844: sine = 32'h4251d5fd;
    11'd845: sine = 32'h4250ca46;
    11'd846: sine = 32'h424fbe0f;
    11'd847: sine = 32'h424eb157;
    11'd848: sine = 32'h424da420;
    11'd849: sine = 32'h424c966a;
    11'd850: sine = 32'h424b8836;
    11'd851: sine = 32'h424a7984;
    11'd852: sine = 32'h42496a56;
    11'd853: sine = 32'h42485aab;
    11'd854: sine = 32'h42474a84;
    11'd855: sine = 32'h424639e3;
    11'd856: sine = 32'h424528c7;
    11'd857: sine = 32'h42441732;
    11'd858: sine = 32'h42430524;
    11'd859: sine = 32'h4241f29d;
    11'd860: sine = 32'h4240df9f;
    11'd861: sine = 32'h423fcc2a;
    11'd862: sine = 32'h423eb83f;
    11'd863: sine = 32'h423da3de;
    11'd864: sine = 32'h423c8f08;
    11'd865: sine = 32'h423b79bd;
    11'd866: sine = 32'h423a63ff;
    11'd867: sine = 32'h42394dce;
    11'd868: sine = 32'h4238372b;
    11'd869: sine = 32'h42372016;
    11'd870: sine = 32'h42360890;
    11'd871: sine = 32'h4234f09a;
    11'd872: sine = 32'h4233d834;
    11'd873: sine = 32'h4232bf60;
    11'd874: sine = 32'h4231a61d;
    11'd875: sine = 32'h42308c6c;
    11'd876: sine = 32'h422f724f;
    11'd877: sine = 32'h422e57c5;
    11'd878: sine = 32'h422d3cd0;
    11'd879: sine = 32'h422c2170;
    11'd880: sine = 32'h422b05a5;
    11'd881: sine = 32'h4229e972;
    11'd882: sine = 32'h4228ccd5;
    11'd883: sine = 32'h4227afd0;
    11'd884: sine = 32'h42269264;
    11'd885: sine = 32'h42257491;
    11'd886: sine = 32'h42245658;
    11'd887: sine = 32'h422337ba;
    11'd888: sine = 32'h422218b7;
    11'd889: sine = 32'h4220f950;
    11'd890: sine = 32'h421fd986;
    11'd891: sine = 32'h421eb959;
    11'd892: sine = 32'h421d98ca;
    11'd893: sine = 32'h421c77da;
    11'd894: sine = 32'h421b568a;
    11'd895: sine = 32'h421a34d9;
    11'd896: sine = 32'h421912ca;
    11'd897: sine = 32'h4217f05c;
    11'd898: sine = 32'h4216cd90;
    11'd899: sine = 32'h4215aa68;
    11'd900: sine = 32'h421486e3;
    11'd901: sine = 32'h42136302;
    11'd902: sine = 32'h42123ec7;
    11'd903: sine = 32'h42111a31;
    11'd904: sine = 32'h420ff542;
    11'd905: sine = 32'h420ecffa;
    11'd906: sine = 32'h420daa59;
    11'd907: sine = 32'h420c8462;
    11'd908: sine = 32'h420b5e14;
    11'd909: sine = 32'h420a3770;
    11'd910: sine = 32'h42091076;
    11'd911: sine = 32'h4207e928;
    11'd912: sine = 32'h4206c187;
    11'd913: sine = 32'h42059992;
    11'd914: sine = 32'h4204714a;
    11'd915: sine = 32'h420348b1;
    11'd916: sine = 32'h42021fc7;
    11'd917: sine = 32'h4200f68d;
    11'd918: sine = 32'h41ff9a06;
    11'd919: sine = 32'h41fd4655;
    11'd920: sine = 32'h41faf208;
    11'd921: sine = 32'h41f89d1f;
    11'd922: sine = 32'h41f6479e;
    11'd923: sine = 32'h41f3f184;
    11'd924: sine = 32'h41f19ad4;
    11'd925: sine = 32'h41ef438f;
    11'd926: sine = 32'h41ecebb6;
    11'd927: sine = 32'h41ea934b;
    11'd928: sine = 32'h41e83a50;
    11'd929: sine = 32'h41e5e0c5;
    11'd930: sine = 32'h41e386ac;
    11'd931: sine = 32'h41e12c07;
    11'd932: sine = 32'h41ded0d8;
    11'd933: sine = 32'h41dc751e;
    11'd934: sine = 32'h41da18dd;
    11'd935: sine = 32'h41d7bc15;
    11'd936: sine = 32'h41d55ec8;
    11'd937: sine = 32'h41d300f8;
    11'd938: sine = 32'h41d0a2a5;
    11'd939: sine = 32'h41ce43d2;
    11'd940: sine = 32'h41cbe47f;
    11'd941: sine = 32'h41c984af;
    11'd942: sine = 32'h41c72462;
    11'd943: sine = 32'h41c4c39b;
    11'd944: sine = 32'h41c2625a;
    11'd945: sine = 32'h41c000a1;
    11'd946: sine = 32'h41bd9e72;
    11'd947: sine = 32'h41bb3bce;
    11'd948: sine = 32'h41b8d8b6;
    11'd949: sine = 32'h41b6752c;
    11'd950: sine = 32'h41b41132;
    11'd951: sine = 32'h41b1acc9;
    11'd952: sine = 32'h41af47f2;
    11'd953: sine = 32'h41ace2af;
    11'd954: sine = 32'h41aa7d01;
    11'd955: sine = 32'h41a816ea;
    11'd956: sine = 32'h41a5b06b;
    11'd957: sine = 32'h41a34987;
    11'd958: sine = 32'h41a0e23d;
    11'd959: sine = 32'h419e7a91;
    11'd960: sine = 32'h419c1282;
    11'd961: sine = 32'h4199aa13;
    11'd962: sine = 32'h41974146;
    11'd963: sine = 32'h4194d81b;
    11'd964: sine = 32'h41926e94;
    11'd965: sine = 32'h419004b3;
    11'd966: sine = 32'h418d9a79;
    11'd967: sine = 32'h418b2fe8;
    11'd968: sine = 32'h4188c501;
    11'd969: sine = 32'h418659c6;
    11'd970: sine = 32'h4183ee38;
    11'd971: sine = 32'h41818258;
    11'd972: sine = 32'h417e2c51;
    11'd973: sine = 32'h41795355;
    11'd974: sine = 32'h417479bf;
    11'd975: sine = 32'h416f9f93;
    11'd976: sine = 32'h416ac4d3;
    11'd977: sine = 32'h4165e982;
    11'd978: sine = 32'h41610da3;
    11'd979: sine = 32'h415c3139;
    11'd980: sine = 32'h41575447;
    11'd981: sine = 32'h415276d1;
    11'd982: sine = 32'h414d98d9;
    11'd983: sine = 32'h4148ba62;
    11'd984: sine = 32'h4143db6f;
    11'd985: sine = 32'h413efc03;
    11'd986: sine = 32'h413a1c22;
    11'd987: sine = 32'h41353bce;
    11'd988: sine = 32'h41305b0a;
    11'd989: sine = 32'h412b79d9;
    11'd990: sine = 32'h4126983e;
    11'd991: sine = 32'h4121b63d;
    11'd992: sine = 32'h411cd3d8;
    11'd993: sine = 32'h4117f112;
    11'd994: sine = 32'h41130dee;
    11'd995: sine = 32'h410e2a70;
    11'd996: sine = 32'h4109469a;
    11'd997: sine = 32'h4104626f;
    11'd998: sine = 32'h40fefbe5;
    11'd999: sine = 32'h40f5324f;
    11'd1000: sine = 32'h40eb6822;
    11'd1001: sine = 32'h40e19d64;
    11'd1002: sine = 32'h40d7d21a;
    11'd1003: sine = 32'h40ce064b;
    11'd1004: sine = 32'h40c439fd;
    11'd1005: sine = 32'h40ba6d37;
    11'd1006: sine = 32'h40b09ffd;
    11'd1007: sine = 32'h40a6d256;
    11'd1008: sine = 32'h409d0448;
    11'd1009: sine = 32'h409335da;
    11'd1010: sine = 32'h40896710;
    11'd1011: sine = 32'h407f2fe4;
    11'd1012: sine = 32'h406b910a;
    11'd1013: sine = 32'h4057f19f;
    11'd1014: sine = 32'h404451af;
    11'd1015: sine = 32'h4030b146;
    11'd1016: sine = 32'h401d1070;
    11'd1017: sine = 32'h40096f38;
    11'd1018: sine = 32'h3feb9b59;
    11'd1019: sine = 32'h3fc457b0;
    11'd1020: sine = 32'h3f9d138d;
    11'd1021: sine = 32'h3f6b9e14;
    11'd1022: sine = 32'h3f1d147c;
    11'd1023: sine = 32'h3e9d1506;
    11'd1024: sine = 32'h36b3d148;
    11'd1025: sine = 32'hbe9d139f;
    11'd1026: sine = 32'hbf1d13c8;
    11'd1027: sine = 32'hbf6b9d60;
    11'd1028: sine = 32'hbf9d1333;
    11'd1029: sine = 32'hbfc45756;
    11'd1030: sine = 32'hbfeb9aff;
    11'd1031: sine = 32'hc0096f0b;
    11'd1032: sine = 32'hc01d1043;
    11'd1033: sine = 32'hc030b119;
    11'd1034: sine = 32'hc0445182;
    11'd1035: sine = 32'hc057f173;
    11'd1036: sine = 32'hc06b90de;
    11'd1037: sine = 32'hc07f2fb7;
    11'd1038: sine = 32'hc08966fa;
    11'd1039: sine = 32'hc09335c3;
    11'd1040: sine = 32'hc09d0432;
    11'd1041: sine = 32'hc0a6d23f;
    11'd1042: sine = 32'hc0b09fe6;
    11'd1043: sine = 32'hc0ba6d20;
    11'd1044: sine = 32'hc0c439e7;
    11'd1045: sine = 32'hc0ce0635;
    11'd1046: sine = 32'hc0d7d204;
    11'd1047: sine = 32'hc0e19d4d;
    11'd1048: sine = 32'hc0eb680c;
    11'd1049: sine = 32'hc0f53239;
    11'd1050: sine = 32'hc0fefbcf;
    11'd1051: sine = 32'hc1046264;
    11'd1052: sine = 32'hc109468f;
    11'd1053: sine = 32'hc10e2a65;
    11'd1054: sine = 32'hc1130de3;
    11'd1055: sine = 32'hc117f106;
    11'd1056: sine = 32'hc11cd3cc;
    11'd1057: sine = 32'hc121b631;
    11'd1058: sine = 32'hc1269833;
    11'd1059: sine = 32'hc12b79cd;
    11'd1060: sine = 32'hc1305afe;
    11'd1061: sine = 32'hc1353bc2;
    11'd1062: sine = 32'hc13a1c17;
    11'd1063: sine = 32'hc13efbf8;
    11'd1064: sine = 32'hc143db64;
    11'd1065: sine = 32'hc148ba57;
    11'd1066: sine = 32'hc14d98ce;
    11'd1067: sine = 32'hc15276c6;
    11'd1068: sine = 32'hc157543c;
    11'd1069: sine = 32'hc15c312e;
    11'd1070: sine = 32'hc1610d98;
    11'd1071: sine = 32'hc165e976;
    11'd1072: sine = 32'hc16ac4c8;
    11'd1073: sine = 32'hc16f9f88;
    11'd1074: sine = 32'hc17479b4;
    11'd1075: sine = 32'hc179534a;
    11'd1076: sine = 32'hc17e2c46;
    11'd1077: sine = 32'hc1818252;
    11'd1078: sine = 32'hc183ee32;
    11'd1079: sine = 32'hc18659c0;
    11'd1080: sine = 32'hc188c4fc;
    11'd1081: sine = 32'hc18b2fe3;
    11'd1082: sine = 32'hc18d9a74;
    11'd1083: sine = 32'hc19004ae;
    11'd1084: sine = 32'hc1926e8f;
    11'd1085: sine = 32'hc194d815;
    11'd1086: sine = 32'hc1974140;
    11'd1087: sine = 32'hc199aa0e;
    11'd1088: sine = 32'hc19c127d;
    11'd1089: sine = 32'hc19e7a8b;
    11'd1090: sine = 32'hc1a0e238;
    11'd1091: sine = 32'hc1a34981;
    11'd1092: sine = 32'hc1a5b066;
    11'd1093: sine = 32'hc1a816e5;
    11'd1094: sine = 32'hc1aa7cfb;
    11'd1095: sine = 32'hc1ace2a9;
    11'd1096: sine = 32'hc1af47ec;
    11'd1097: sine = 32'hc1b1acc3;
    11'd1098: sine = 32'hc1b4112c;
    11'd1099: sine = 32'hc1b67527;
    11'd1100: sine = 32'hc1b8d8b0;
    11'd1101: sine = 32'hc1bb3bc8;
    11'd1102: sine = 32'hc1bd9e6c;
    11'd1103: sine = 32'hc1c0009c;
    11'd1104: sine = 32'hc1c26254;
    11'd1105: sine = 32'hc1c4c395;
    11'd1106: sine = 32'hc1c7245d;
    11'd1107: sine = 32'hc1c984a9;
    11'd1108: sine = 32'hc1cbe47a;
    11'd1109: sine = 32'hc1ce43cc;
    11'd1110: sine = 32'hc1d0a2a0;
    11'd1111: sine = 32'hc1d300f2;
    11'd1112: sine = 32'hc1d55ec3;
    11'd1113: sine = 32'hc1d7bc10;
    11'd1114: sine = 32'hc1da18d8;
    11'd1115: sine = 32'hc1dc7519;
    11'd1116: sine = 32'hc1ded0d2;
    11'd1117: sine = 32'hc1e12c02;
    11'd1118: sine = 32'hc1e386a7;
    11'd1119: sine = 32'hc1e5e0c0;
    11'd1120: sine = 32'hc1e83a4a;
    11'd1121: sine = 32'hc1ea9346;
    11'd1122: sine = 32'hc1ecebb1;
    11'd1123: sine = 32'hc1ef4389;
    11'd1124: sine = 32'hc1f19acf;
    11'd1125: sine = 32'hc1f3f17f;
    11'd1126: sine = 32'hc1f64798;
    11'd1127: sine = 32'hc1f89d1a;
    11'd1128: sine = 32'hc1faf202;
    11'd1129: sine = 32'hc1fd4650;
    11'd1130: sine = 32'hc1ff9a01;
    11'd1131: sine = 32'hc200f68a;
    11'd1132: sine = 32'hc2021fc5;
    11'd1133: sine = 32'hc20348af;
    11'd1134: sine = 32'hc2047148;
    11'd1135: sine = 32'hc205998f;
    11'd1136: sine = 32'hc206c184;
    11'd1137: sine = 32'hc207e926;
    11'd1138: sine = 32'hc2091074;
    11'd1139: sine = 32'hc20a376d;
    11'd1140: sine = 32'hc20b5e11;
    11'd1141: sine = 32'hc20c845f;
    11'd1142: sine = 32'hc20daa57;
    11'd1143: sine = 32'hc20ecff7;
    11'd1144: sine = 32'hc20ff53f;
    11'd1145: sine = 32'hc2111a2e;
    11'd1146: sine = 32'hc2123ec4;
    11'd1147: sine = 32'hc21362ff;
    11'd1148: sine = 32'hc21486e0;
    11'd1149: sine = 32'hc215aa65;
    11'd1150: sine = 32'hc216cd8e;
    11'd1151: sine = 32'hc217f059;
    11'd1152: sine = 32'hc21912c7;
    11'd1153: sine = 32'hc21a34d7;
    11'd1154: sine = 32'hc21b5687;
    11'd1155: sine = 32'hc21c77d7;
    11'd1156: sine = 32'hc21d98c7;
    11'd1157: sine = 32'hc21eb956;
    11'd1158: sine = 32'hc21fd983;
    11'd1159: sine = 32'hc220f94d;
    11'd1160: sine = 32'hc22218b4;
    11'd1161: sine = 32'hc22337b7;
    11'd1162: sine = 32'hc2245656;
    11'd1163: sine = 32'hc225748f;
    11'd1164: sine = 32'hc2269262;
    11'd1165: sine = 32'hc227afce;
    11'd1166: sine = 32'hc228ccd2;
    11'd1167: sine = 32'hc229e96f;
    11'd1168: sine = 32'hc22b05a3;
    11'd1169: sine = 32'hc22c216d;
    11'd1170: sine = 32'hc22d3ccd;
    11'd1171: sine = 32'hc22e57c2;
    11'd1172: sine = 32'hc22f724c;
    11'd1173: sine = 32'hc2308c6a;
    11'd1174: sine = 32'hc231a61a;
    11'd1175: sine = 32'hc232bf5d;
    11'd1176: sine = 32'hc233d832;
    11'd1177: sine = 32'hc234f098;
    11'd1178: sine = 32'hc236088e;
    11'd1179: sine = 32'hc2372014;
    11'd1180: sine = 32'hc2383729;
    11'd1181: sine = 32'hc2394dcc;
    11'd1182: sine = 32'hc23a63fd;
    11'd1183: sine = 32'hc23b79bb;
    11'd1184: sine = 32'hc23c8f05;
    11'd1185: sine = 32'hc23da3db;
    11'd1186: sine = 32'hc23eb83c;
    11'd1187: sine = 32'hc23fcc28;
    11'd1188: sine = 32'hc240df9d;
    11'd1189: sine = 32'hc241f29b;
    11'd1190: sine = 32'hc2430521;
    11'd1191: sine = 32'hc2441730;
    11'd1192: sine = 32'hc24528c5;
    11'd1193: sine = 32'hc24639e1;
    11'd1194: sine = 32'hc2474a82;
    11'd1195: sine = 32'hc2485aa8;
    11'd1196: sine = 32'hc2496a53;
    11'd1197: sine = 32'hc24a7982;
    11'd1198: sine = 32'hc24b8833;
    11'd1199: sine = 32'hc24c9668;
    11'd1200: sine = 32'hc24da41e;
    11'd1201: sine = 32'hc24eb155;
    11'd1202: sine = 32'hc24fbe0c;
    11'd1203: sine = 32'hc250ca44;
    11'd1204: sine = 32'hc251d5fa;
    11'd1205: sine = 32'hc252e130;
    11'd1206: sine = 32'hc253ebe3;
    11'd1207: sine = 32'hc254f613;
    11'd1208: sine = 32'hc255ffc0;
    11'd1209: sine = 32'hc25708e9;
    11'd1210: sine = 32'hc258118e;
    11'd1211: sine = 32'hc25919ad;
    11'd1212: sine = 32'hc25a2146;
    11'd1213: sine = 32'hc25b2859;
    11'd1214: sine = 32'hc25c2ee4;
    11'd1215: sine = 32'hc25d34e8;
    11'd1216: sine = 32'hc25e3a63;
    11'd1217: sine = 32'hc25f3f55;
    11'd1218: sine = 32'hc26043bd;
    11'd1219: sine = 32'hc261479c;
    11'd1220: sine = 32'hc2624aef;
    11'd1221: sine = 32'hc2634db6;
    11'd1222: sine = 32'hc2644ff1;
    11'd1223: sine = 32'hc26551a0;
    11'd1224: sine = 32'hc26652c1;
    11'd1225: sine = 32'hc2675354;
    11'd1226: sine = 32'hc2685358;
    11'd1227: sine = 32'hc26952cd;
    11'd1228: sine = 32'hc26a51b2;
    11'd1229: sine = 32'hc26b5006;
    11'd1230: sine = 32'hc26c4dca;
    11'd1231: sine = 32'hc26d4afb;
    11'd1232: sine = 32'hc26e479a;
    11'd1233: sine = 32'hc26f43a7;
    11'd1234: sine = 32'hc2703f1f;
    11'd1235: sine = 32'hc2713a04;
    11'd1236: sine = 32'hc2723453;
    11'd1237: sine = 32'hc2732e0d;
    11'd1238: sine = 32'hc2742732;
    11'd1239: sine = 32'hc2751fbf;
    11'd1240: sine = 32'hc27617b6;
    11'd1241: sine = 32'hc2770f14;
    11'd1242: sine = 32'hc27805da;
    11'd1243: sine = 32'hc278fc08;
    11'd1244: sine = 32'hc279f19b;
    11'd1245: sine = 32'hc27ae695;
    11'd1246: sine = 32'hc27bdaf3;
    11'd1247: sine = 32'hc27cceb7;
    11'd1248: sine = 32'hc27dc1de;
    11'd1249: sine = 32'hc27eb469;
    11'd1250: sine = 32'hc27fa657;
    11'd1251: sine = 32'hc2804bd3;
    11'd1252: sine = 32'hc280c42c;
    11'd1253: sine = 32'hc2813c36;
    11'd1254: sine = 32'hc281b3ef;
    11'd1255: sine = 32'hc2822b59;
    11'd1256: sine = 32'hc282a272;
    11'd1257: sine = 32'hc283193b;
    11'd1258: sine = 32'hc2838fb3;
    11'd1259: sine = 32'hc28405da;
    11'd1260: sine = 32'hc2847baf;
    11'd1261: sine = 32'hc284f133;
    11'd1262: sine = 32'hc2856665;
    11'd1263: sine = 32'hc285db44;
    11'd1264: sine = 32'hc2864fd1;
    11'd1265: sine = 32'hc286c40b;
    11'd1266: sine = 32'hc28737f2;
    11'd1267: sine = 32'hc287ab85;
    11'd1268: sine = 32'hc2881ec5;
    11'd1269: sine = 32'hc28891b1;
    11'd1270: sine = 32'hc2890448;
    11'd1271: sine = 32'hc289768b;
    11'd1272: sine = 32'hc289e879;
    11'd1273: sine = 32'hc28a5a12;
    11'd1274: sine = 32'hc28acb56;
    11'd1275: sine = 32'hc28b3c44;
    11'd1276: sine = 32'hc28bacdd;
    11'd1277: sine = 32'hc28c1d1f;
    11'd1278: sine = 32'hc28c8d0a;
    11'd1279: sine = 32'hc28cfc9f;
    11'd1280: sine = 32'hc28d6bdd;
    11'd1281: sine = 32'hc28ddac4;
    11'd1282: sine = 32'hc28e4953;
    11'd1283: sine = 32'hc28eb78b;
    11'd1284: sine = 32'hc28f256a;
    11'd1285: sine = 32'hc28f92f2;
    11'd1286: sine = 32'hc2900020;
    11'd1287: sine = 32'hc2906cf6;
    11'd1288: sine = 32'hc290d973;
    11'd1289: sine = 32'hc2914596;
    11'd1290: sine = 32'hc291b160;
    11'd1291: sine = 32'hc2921cd0;
    11'd1292: sine = 32'hc29287e5;
    11'd1293: sine = 32'hc292f2a1;
    11'd1294: sine = 32'hc2935d02;
    11'd1295: sine = 32'hc293c707;
    11'd1296: sine = 32'hc29430b2;
    11'd1297: sine = 32'hc2949a01;
    11'd1298: sine = 32'hc29502f5;
    11'd1299: sine = 32'hc2956b8c;
    11'd1300: sine = 32'hc295d3c8;
    11'd1301: sine = 32'hc2963ba7;
    11'd1302: sine = 32'hc296a329;
    11'd1303: sine = 32'hc2970a4f;
    11'd1304: sine = 32'hc2977117;
    11'd1305: sine = 32'hc297d782;
    11'd1306: sine = 32'hc2983d8f;
    11'd1307: sine = 32'hc298a33f;
    11'd1308: sine = 32'hc2990890;
    11'd1309: sine = 32'hc2996d83;
    11'd1310: sine = 32'hc299d217;
    11'd1311: sine = 32'hc29a364c;
    11'd1312: sine = 32'hc29a9a22;
    11'd1313: sine = 32'hc29afd99;
    11'd1314: sine = 32'hc29b60b0;
    11'd1315: sine = 32'hc29bc367;
    11'd1316: sine = 32'hc29c25be;
    11'd1317: sine = 32'hc29c87b5;
    11'd1318: sine = 32'hc29ce94c;
    11'd1319: sine = 32'hc29d4a81;
    11'd1320: sine = 32'hc29dab56;
    11'd1321: sine = 32'hc29e0bc9;
    11'd1322: sine = 32'hc29e6bdb;
    11'd1323: sine = 32'hc29ecb8b;
    11'd1324: sine = 32'hc29f2ad9;
    11'd1325: sine = 32'hc29f89c5;
    11'd1326: sine = 32'hc29fe84e;
    11'd1327: sine = 32'hc2a04675;
    11'd1328: sine = 32'hc2a0a439;
    11'd1329: sine = 32'hc2a1019a;
    11'd1330: sine = 32'hc2a15e98;
    11'd1331: sine = 32'hc2a1bb32;
    11'd1332: sine = 32'hc2a21768;
    11'd1333: sine = 32'hc2a2733a;
    11'd1334: sine = 32'hc2a2cea8;
    11'd1335: sine = 32'hc2a329b2;
    11'd1336: sine = 32'hc2a38457;
    11'd1337: sine = 32'hc2a3de97;
    11'd1338: sine = 32'hc2a43872;
    11'd1339: sine = 32'hc2a491e8;
    11'd1340: sine = 32'hc2a4eaf8;
    11'd1341: sine = 32'hc2a543a3;
    11'd1342: sine = 32'hc2a59be8;
    11'd1343: sine = 32'hc2a5f3c6;
    11'd1344: sine = 32'hc2a64b3e;
    11'd1345: sine = 32'hc2a6a24f;
    11'd1346: sine = 32'hc2a6f8fa;
    11'd1347: sine = 32'hc2a74f3e;
    11'd1348: sine = 32'hc2a7a51a;
    11'd1349: sine = 32'hc2a7fa8f;
    11'd1350: sine = 32'hc2a84f9d;
    11'd1351: sine = 32'hc2a8a443;
    11'd1352: sine = 32'hc2a8f880;
    11'd1353: sine = 32'hc2a94c56;
    11'd1354: sine = 32'hc2a99fc2;
    11'd1355: sine = 32'hc2a9f2c7;
    11'd1356: sine = 32'hc2aa4562;
    11'd1357: sine = 32'hc2aa9795;
    11'd1358: sine = 32'hc2aae95e;
    11'd1359: sine = 32'hc2ab3abe;
    11'd1360: sine = 32'hc2ab8bb4;
    11'd1361: sine = 32'hc2abdc40;
    11'd1362: sine = 32'hc2ac2c63;
    11'd1363: sine = 32'hc2ac7c1b;
    11'd1364: sine = 32'hc2accb69;
    11'd1365: sine = 32'hc2ad1a4c;
    11'd1366: sine = 32'hc2ad68c4;
    11'd1367: sine = 32'hc2adb6d1;
    11'd1368: sine = 32'hc2ae0474;
    11'd1369: sine = 32'hc2ae51ab;
    11'd1370: sine = 32'hc2ae9e76;
    11'd1371: sine = 32'hc2aeead6;
    11'd1372: sine = 32'hc2af36c9;
    11'd1373: sine = 32'hc2af8251;
    11'd1374: sine = 32'hc2afcd6d;
    11'd1375: sine = 32'hc2b0181c;
    11'd1376: sine = 32'hc2b0625e;
    11'd1377: sine = 32'hc2b0ac34;
    11'd1378: sine = 32'hc2b0f59c;
    11'd1379: sine = 32'hc2b13e98;
    11'd1380: sine = 32'hc2b18726;
    11'd1381: sine = 32'hc2b1cf46;
    11'd1382: sine = 32'hc2b216f9;
    11'd1383: sine = 32'hc2b25e3e;
    11'd1384: sine = 32'hc2b2a515;
    11'd1385: sine = 32'hc2b2eb7e;
    11'd1386: sine = 32'hc2b33178;
    11'd1387: sine = 32'hc2b37704;
    11'd1388: sine = 32'hc2b3bc22;
    11'd1389: sine = 32'hc2b400d0;
    11'd1390: sine = 32'hc2b4450f;
    11'd1391: sine = 32'hc2b488df;
    11'd1392: sine = 32'hc2b4cc40;
    11'd1393: sine = 32'hc2b50f31;
    11'd1394: sine = 32'hc2b551b3;
    11'd1395: sine = 32'hc2b593c5;
    11'd1396: sine = 32'hc2b5d566;
    11'd1397: sine = 32'hc2b61698;
    11'd1398: sine = 32'hc2b65759;
    11'd1399: sine = 32'hc2b697aa;
    11'd1400: sine = 32'hc2b6d78a;
    11'd1401: sine = 32'hc2b716f9;
    11'd1402: sine = 32'hc2b755f7;
    11'd1403: sine = 32'hc2b79485;
    11'd1404: sine = 32'hc2b7d2a1;
    11'd1405: sine = 32'hc2b8104b;
    11'd1406: sine = 32'hc2b84d84;
    11'd1407: sine = 32'hc2b88a4c;
    11'd1408: sine = 32'hc2b8c6a1;
    11'd1409: sine = 32'hc2b90285;
    11'd1410: sine = 32'hc2b93df7;
    11'd1411: sine = 32'hc2b978f6;
    11'd1412: sine = 32'hc2b9b383;
    11'd1413: sine = 32'hc2b9ed9d;
    11'd1414: sine = 32'hc2ba2744;
    11'd1415: sine = 32'hc2ba6079;
    11'd1416: sine = 32'hc2ba993b;
    11'd1417: sine = 32'hc2bad18a;
    11'd1418: sine = 32'hc2bb0965;
    11'd1419: sine = 32'hc2bb40cd;
    11'd1420: sine = 32'hc2bb77c2;
    11'd1421: sine = 32'hc2bbae42;
    11'd1422: sine = 32'hc2bbe450;
    11'd1423: sine = 32'hc2bc19e9;
    11'd1424: sine = 32'hc2bc4f0e;
    11'd1425: sine = 32'hc2bc83bf;
    11'd1426: sine = 32'hc2bcb7fc;
    11'd1427: sine = 32'hc2bcebc4;
    11'd1428: sine = 32'hc2bd1f18;
    11'd1429: sine = 32'hc2bd51f7;
    11'd1430: sine = 32'hc2bd8462;
    11'd1431: sine = 32'hc2bdb657;
    11'd1432: sine = 32'hc2bde7d7;
    11'd1433: sine = 32'hc2be18e3;
    11'd1434: sine = 32'hc2be4979;
    11'd1435: sine = 32'hc2be7999;
    11'd1436: sine = 32'hc2bea945;
    11'd1437: sine = 32'hc2bed87a;
    11'd1438: sine = 32'hc2bf073a;
    11'd1439: sine = 32'hc2bf3584;
    11'd1440: sine = 32'hc2bf6358;
    11'd1441: sine = 32'hc2bf90b6;
    11'd1442: sine = 32'hc2bfbd9e;
    11'd1443: sine = 32'hc2bfea0f;
    11'd1444: sine = 32'hc2c0160b;
    11'd1445: sine = 32'hc2c0418f;
    11'd1446: sine = 32'hc2c06c9d;
    11'd1447: sine = 32'hc2c09735;
    11'd1448: sine = 32'hc2c0c155;
    11'd1449: sine = 32'hc2c0eaff;
    11'd1450: sine = 32'hc2c11432;
    11'd1451: sine = 32'hc2c13ced;
    11'd1452: sine = 32'hc2c16532;
    11'd1453: sine = 32'hc2c18cff;
    11'd1454: sine = 32'hc2c1b455;
    11'd1455: sine = 32'hc2c1db33;
    11'd1456: sine = 32'hc2c20199;
    11'd1457: sine = 32'hc2c22788;
    11'd1458: sine = 32'hc2c24d00;
    11'd1459: sine = 32'hc2c271ff;
    11'd1460: sine = 32'hc2c29686;
    11'd1461: sine = 32'hc2c2ba96;
    11'd1462: sine = 32'hc2c2de2d;
    11'd1463: sine = 32'hc2c3014c;
    11'd1464: sine = 32'hc2c323f3;
    11'd1465: sine = 32'hc2c34621;
    11'd1466: sine = 32'hc2c367d7;
    11'd1467: sine = 32'hc2c38914;
    11'd1468: sine = 32'hc2c3a9d9;
    11'd1469: sine = 32'hc2c3ca25;
    11'd1470: sine = 32'hc2c3e9f9;
    11'd1471: sine = 32'hc2c40953;
    11'd1472: sine = 32'hc2c42835;
    11'd1473: sine = 32'hc2c4469d;
    11'd1474: sine = 32'hc2c4648d;
    11'd1475: sine = 32'hc2c48203;
    11'd1476: sine = 32'hc2c49f00;
    11'd1477: sine = 32'hc2c4bb84;
    11'd1478: sine = 32'hc2c4d78e;
    11'd1479: sine = 32'hc2c4f31f;
    11'd1480: sine = 32'hc2c50e37;
    11'd1481: sine = 32'hc2c528d5;
    11'd1482: sine = 32'hc2c542f9;
    11'd1483: sine = 32'hc2c55ca4;
    11'd1484: sine = 32'hc2c575d5;
    11'd1485: sine = 32'hc2c58e8c;
    11'd1486: sine = 32'hc2c5a6c9;
    11'd1487: sine = 32'hc2c5be8d;
    11'd1488: sine = 32'hc2c5d5d6;
    11'd1489: sine = 32'hc2c5eca6;
    11'd1490: sine = 32'hc2c602fb;
    11'd1491: sine = 32'hc2c618d6;
    11'd1492: sine = 32'hc2c62e37;
    11'd1493: sine = 32'hc2c6431e;
    11'd1494: sine = 32'hc2c6578a;
    11'd1495: sine = 32'hc2c66b7c;
    11'd1496: sine = 32'hc2c67ef4;
    11'd1497: sine = 32'hc2c691f1;
    11'd1498: sine = 32'hc2c6a474;
    11'd1499: sine = 32'hc2c6b67c;
    11'd1500: sine = 32'hc2c6c809;
    11'd1501: sine = 32'hc2c6d91c;
    11'd1502: sine = 32'hc2c6e9b5;
    11'd1503: sine = 32'hc2c6f9d2;
    11'd1504: sine = 32'hc2c70975;
    11'd1505: sine = 32'hc2c7189d;
    11'd1506: sine = 32'hc2c7274b;
    11'd1507: sine = 32'hc2c7357d;
    11'd1508: sine = 32'hc2c74335;
    11'd1509: sine = 32'hc2c75071;
    11'd1510: sine = 32'hc2c75d33;
    11'd1511: sine = 32'hc2c7697a;
    11'd1512: sine = 32'hc2c77545;
    11'd1513: sine = 32'hc2c78096;
    11'd1514: sine = 32'hc2c78b6c;
    11'd1515: sine = 32'hc2c795c6;
    11'd1516: sine = 32'hc2c79fa6;
    11'd1517: sine = 32'hc2c7a90a;
    11'd1518: sine = 32'hc2c7b1f3;
    11'd1519: sine = 32'hc2c7ba61;
    11'd1520: sine = 32'hc2c7c254;
    11'd1521: sine = 32'hc2c7c9cb;
    11'd1522: sine = 32'hc2c7d0c8;
    11'd1523: sine = 32'hc2c7d749;
    11'd1524: sine = 32'hc2c7dd4e;
    11'd1525: sine = 32'hc2c7e2d9;
    11'd1526: sine = 32'hc2c7e7e8;
    11'd1527: sine = 32'hc2c7ec7c;
    11'd1528: sine = 32'hc2c7f094;
    11'd1529: sine = 32'hc2c7f432;
    11'd1530: sine = 32'hc2c7f753;
    11'd1531: sine = 32'hc2c7f9fa;
    11'd1532: sine = 32'hc2c7fc25;
    11'd1533: sine = 32'hc2c7fdd5;
    11'd1534: sine = 32'hc2c7ff09;
    11'd1535: sine = 32'hc2c7ffc2;
    11'd1536: sine = 32'hc2c80000;
    11'd1537: sine = 32'hc2c7ffc2;
    11'd1538: sine = 32'hc2c7ff09;
    11'd1539: sine = 32'hc2c7fdd5;
    11'd1540: sine = 32'hc2c7fc25;
    11'd1541: sine = 32'hc2c7f9fa;
    11'd1542: sine = 32'hc2c7f753;
    11'd1543: sine = 32'hc2c7f432;
    11'd1544: sine = 32'hc2c7f094;
    11'd1545: sine = 32'hc2c7ec7c;
    11'd1546: sine = 32'hc2c7e7e8;
    11'd1547: sine = 32'hc2c7e2d9;
    11'd1548: sine = 32'hc2c7dd4e;
    11'd1549: sine = 32'hc2c7d749;
    11'd1550: sine = 32'hc2c7d0c8;
    11'd1551: sine = 32'hc2c7c9cb;
    11'd1552: sine = 32'hc2c7c254;
    11'd1553: sine = 32'hc2c7ba61;
    11'd1554: sine = 32'hc2c7b1f3;
    11'd1555: sine = 32'hc2c7a90a;
    11'd1556: sine = 32'hc2c79fa6;
    11'd1557: sine = 32'hc2c795c6;
    11'd1558: sine = 32'hc2c78b6c;
    11'd1559: sine = 32'hc2c78096;
    11'd1560: sine = 32'hc2c77546;
    11'd1561: sine = 32'hc2c7697a;
    11'd1562: sine = 32'hc2c75d33;
    11'd1563: sine = 32'hc2c75071;
    11'd1564: sine = 32'hc2c74335;
    11'd1565: sine = 32'hc2c7357d;
    11'd1566: sine = 32'hc2c7274b;
    11'd1567: sine = 32'hc2c7189d;
    11'd1568: sine = 32'hc2c70975;
    11'd1569: sine = 32'hc2c6f9d2;
    11'd1570: sine = 32'hc2c6e9b5;
    11'd1571: sine = 32'hc2c6d91d;
    11'd1572: sine = 32'hc2c6c80a;
    11'd1573: sine = 32'hc2c6b67c;
    11'd1574: sine = 32'hc2c6a474;
    11'd1575: sine = 32'hc2c691f1;
    11'd1576: sine = 32'hc2c67ef4;
    11'd1577: sine = 32'hc2c66b7c;
    11'd1578: sine = 32'hc2c6578a;
    11'd1579: sine = 32'hc2c6431e;
    11'd1580: sine = 32'hc2c62e37;
    11'd1581: sine = 32'hc2c618d6;
    11'd1582: sine = 32'hc2c602fb;
    11'd1583: sine = 32'hc2c5eca6;
    11'd1584: sine = 32'hc2c5d5d7;
    11'd1585: sine = 32'hc2c5be8d;
    11'd1586: sine = 32'hc2c5a6ca;
    11'd1587: sine = 32'hc2c58e8c;
    11'd1588: sine = 32'hc2c575d5;
    11'd1589: sine = 32'hc2c55ca4;
    11'd1590: sine = 32'hc2c542fa;
    11'd1591: sine = 32'hc2c528d5;
    11'd1592: sine = 32'hc2c50e37;
    11'd1593: sine = 32'hc2c4f320;
    11'd1594: sine = 32'hc2c4d78f;
    11'd1595: sine = 32'hc2c4bb84;
    11'd1596: sine = 32'hc2c49f00;
    11'd1597: sine = 32'hc2c48203;
    11'd1598: sine = 32'hc2c4648d;
    11'd1599: sine = 32'hc2c4469e;
    11'd1600: sine = 32'hc2c42835;
    11'd1601: sine = 32'hc2c40954;
    11'd1602: sine = 32'hc2c3e9f9;
    11'd1603: sine = 32'hc2c3ca26;
    11'd1604: sine = 32'hc2c3a9da;
    11'd1605: sine = 32'hc2c38915;
    11'd1606: sine = 32'hc2c367d8;
    11'd1607: sine = 32'hc2c34622;
    11'd1608: sine = 32'hc2c323f3;
    11'd1609: sine = 32'hc2c3014c;
    11'd1610: sine = 32'hc2c2de2d;
    11'd1611: sine = 32'hc2c2ba96;
    11'd1612: sine = 32'hc2c29687;
    11'd1613: sine = 32'hc2c271ff;
    11'd1614: sine = 32'hc2c24d00;
    11'd1615: sine = 32'hc2c22789;
    11'd1616: sine = 32'hc2c2019a;
    11'd1617: sine = 32'hc2c1db33;
    11'd1618: sine = 32'hc2c1b455;
    11'd1619: sine = 32'hc2c18cff;
    11'd1620: sine = 32'hc2c16532;
    11'd1621: sine = 32'hc2c13cee;
    11'd1622: sine = 32'hc2c11432;
    11'd1623: sine = 32'hc2c0eb00;
    11'd1624: sine = 32'hc2c0c156;
    11'd1625: sine = 32'hc2c09735;
    11'd1626: sine = 32'hc2c06c9e;
    11'd1627: sine = 32'hc2c04190;
    11'd1628: sine = 32'hc2c0160b;
    11'd1629: sine = 32'hc2bfea10;
    11'd1630: sine = 32'hc2bfbd9f;
    11'd1631: sine = 32'hc2bf90b7;
    11'd1632: sine = 32'hc2bf6359;
    11'd1633: sine = 32'hc2bf3585;
    11'd1634: sine = 32'hc2bf073b;
    11'd1635: sine = 32'hc2bed87b;
    11'd1636: sine = 32'hc2bea945;
    11'd1637: sine = 32'hc2be799a;
    11'd1638: sine = 32'hc2be4979;
    11'd1639: sine = 32'hc2be18e3;
    11'd1640: sine = 32'hc2bde7d8;
    11'd1641: sine = 32'hc2bdb658;
    11'd1642: sine = 32'hc2bd8462;
    11'd1643: sine = 32'hc2bd51f8;
    11'd1644: sine = 32'hc2bd1f19;
    11'd1645: sine = 32'hc2bcebc5;
    11'd1646: sine = 32'hc2bcb7fd;
    11'd1647: sine = 32'hc2bc83c0;
    11'd1648: sine = 32'hc2bc4f0f;
    11'd1649: sine = 32'hc2bc19ea;
    11'd1650: sine = 32'hc2bbe450;
    11'd1651: sine = 32'hc2bbae43;
    11'd1652: sine = 32'hc2bb77c2;
    11'd1653: sine = 32'hc2bb40ce;
    11'd1654: sine = 32'hc2bb0966;
    11'd1655: sine = 32'hc2bad18a;
    11'd1656: sine = 32'hc2ba993c;
    11'd1657: sine = 32'hc2ba607a;
    11'd1658: sine = 32'hc2ba2745;
    11'd1659: sine = 32'hc2b9ed9e;
    11'd1660: sine = 32'hc2b9b383;
    11'd1661: sine = 32'hc2b978f7;
    11'd1662: sine = 32'hc2b93df7;
    11'd1663: sine = 32'hc2b90286;
    11'd1664: sine = 32'hc2b8c6a2;
    11'd1665: sine = 32'hc2b88a4d;
    11'd1666: sine = 32'hc2b84d85;
    11'd1667: sine = 32'hc2b8104c;
    11'd1668: sine = 32'hc2b7d2a2;
    11'd1669: sine = 32'hc2b79486;
    11'd1670: sine = 32'hc2b755f8;
    11'd1671: sine = 32'hc2b716fa;
    11'd1672: sine = 32'hc2b6d78b;
    11'd1673: sine = 32'hc2b697aa;
    11'd1674: sine = 32'hc2b6575a;
    11'd1675: sine = 32'hc2b61699;
    11'd1676: sine = 32'hc2b5d567;
    11'd1677: sine = 32'hc2b593c5;
    11'd1678: sine = 32'hc2b551b4;
    11'd1679: sine = 32'hc2b50f32;
    11'd1680: sine = 32'hc2b4cc41;
    11'd1681: sine = 32'hc2b488e0;
    11'd1682: sine = 32'hc2b44510;
    11'd1683: sine = 32'hc2b400d1;
    11'd1684: sine = 32'hc2b3bc22;
    11'd1685: sine = 32'hc2b37705;
    11'd1686: sine = 32'hc2b33179;
    11'd1687: sine = 32'hc2b2eb7f;
    11'd1688: sine = 32'hc2b2a516;
    11'd1689: sine = 32'hc2b25e3f;
    11'd1690: sine = 32'hc2b216fa;
    11'd1691: sine = 32'hc2b1cf47;
    11'd1692: sine = 32'hc2b18727;
    11'd1693: sine = 32'hc2b13e98;
    11'd1694: sine = 32'hc2b0f59d;
    11'd1695: sine = 32'hc2b0ac34;
    11'd1696: sine = 32'hc2b0625f;
    11'd1697: sine = 32'hc2b0181d;
    11'd1698: sine = 32'hc2afcd6e;
    11'd1699: sine = 32'hc2af8252;
    11'd1700: sine = 32'hc2af36cb;
    11'd1701: sine = 32'hc2aeead7;
    11'd1702: sine = 32'hc2ae9e77;
    11'd1703: sine = 32'hc2ae51ac;
    11'd1704: sine = 32'hc2ae0475;
    11'd1705: sine = 32'hc2adb6d3;
    11'd1706: sine = 32'hc2ad68c5;
    11'd1707: sine = 32'hc2ad1a4d;
    11'd1708: sine = 32'hc2accb6a;
    11'd1709: sine = 32'hc2ac7c1c;
    11'd1710: sine = 32'hc2ac2c64;
    11'd1711: sine = 32'hc2abdc41;
    11'd1712: sine = 32'hc2ab8bb5;
    11'd1713: sine = 32'hc2ab3abf;
    11'd1714: sine = 32'hc2aae95f;
    11'd1715: sine = 32'hc2aa9796;
    11'd1716: sine = 32'hc2aa4563;
    11'd1717: sine = 32'hc2a9f2c8;
    11'd1718: sine = 32'hc2a99fc4;
    11'd1719: sine = 32'hc2a94c57;
    11'd1720: sine = 32'hc2a8f881;
    11'd1721: sine = 32'hc2a8a444;
    11'd1722: sine = 32'hc2a84f9e;
    11'd1723: sine = 32'hc2a7fa91;
    11'd1724: sine = 32'hc2a7a51c;
    11'd1725: sine = 32'hc2a74f3f;
    11'd1726: sine = 32'hc2a6f8fb;
    11'd1727: sine = 32'hc2a6a251;
    11'd1728: sine = 32'hc2a64b3f;
    11'd1729: sine = 32'hc2a5f3c7;
    11'd1730: sine = 32'hc2a59be9;
    11'd1731: sine = 32'hc2a543a4;
    11'd1732: sine = 32'hc2a4eafa;
    11'd1733: sine = 32'hc2a491e9;
    11'd1734: sine = 32'hc2a43874;
    11'd1735: sine = 32'hc2a3de98;
    11'd1736: sine = 32'hc2a38458;
    11'd1737: sine = 32'hc2a329b3;
    11'd1738: sine = 32'hc2a2ceaa;
    11'd1739: sine = 32'hc2a2733c;
    11'd1740: sine = 32'hc2a21769;
    11'd1741: sine = 32'hc2a1bb33;
    11'd1742: sine = 32'hc2a15e99;
    11'd1743: sine = 32'hc2a1019b;
    11'd1744: sine = 32'hc2a0a43a;
    11'd1745: sine = 32'hc2a04676;
    11'd1746: sine = 32'hc29fe850;
    11'd1747: sine = 32'hc29f89c6;
    11'd1748: sine = 32'hc29f2ada;
    11'd1749: sine = 32'hc29ecb8c;
    11'd1750: sine = 32'hc29e6bdc;
    11'd1751: sine = 32'hc29e0bca;
    11'd1752: sine = 32'hc29dab57;
    11'd1753: sine = 32'hc29d4a83;
    11'd1754: sine = 32'hc29ce94d;
    11'd1755: sine = 32'hc29c87b7;
    11'd1756: sine = 32'hc29c25c0;
    11'd1757: sine = 32'hc29bc369;
    11'd1758: sine = 32'hc29b60b1;
    11'd1759: sine = 32'hc29afd9a;
    11'd1760: sine = 32'hc29a9a23;
    11'd1761: sine = 32'hc29a364d;
    11'd1762: sine = 32'hc299d218;
    11'd1763: sine = 32'hc2996d84;
    11'd1764: sine = 32'hc2990891;
    11'd1765: sine = 32'hc298a340;
    11'd1766: sine = 32'hc2983d91;
    11'd1767: sine = 32'hc297d783;
    11'd1768: sine = 32'hc2977119;
    11'd1769: sine = 32'hc2970a50;
    11'd1770: sine = 32'hc296a32b;
    11'd1771: sine = 32'hc2963ba8;
    11'd1772: sine = 32'hc295d3c9;
    11'd1773: sine = 32'hc2956b8e;
    11'd1774: sine = 32'hc29502f6;
    11'd1775: sine = 32'hc2949a03;
    11'd1776: sine = 32'hc29430b3;
    11'd1777: sine = 32'hc293c709;
    11'd1778: sine = 32'hc2935d03;
    11'd1779: sine = 32'hc292f2a2;
    11'd1780: sine = 32'hc29287e7;
    11'd1781: sine = 32'hc2921cd1;
    11'd1782: sine = 32'hc291b161;
    11'd1783: sine = 32'hc2914598;
    11'd1784: sine = 32'hc290d974;
    11'd1785: sine = 32'hc2906cf8;
    11'd1786: sine = 32'hc2900022;
    11'd1787: sine = 32'hc28f92f3;
    11'd1788: sine = 32'hc28f256c;
    11'd1789: sine = 32'hc28eb78c;
    11'd1790: sine = 32'hc28e4955;
    11'd1791: sine = 32'hc28ddac6;
    11'd1792: sine = 32'hc28d6bdf;
    11'd1793: sine = 32'hc28cfca1;
    11'd1794: sine = 32'hc28c8d0c;
    11'd1795: sine = 32'hc28c1d20;
    11'd1796: sine = 32'hc28bacde;
    11'd1797: sine = 32'hc28b3c46;
    11'd1798: sine = 32'hc28acb58;
    11'd1799: sine = 32'hc28a5a14;
    11'd1800: sine = 32'hc289e87b;
    11'd1801: sine = 32'hc289768d;
    11'd1802: sine = 32'hc289044a;
    11'd1803: sine = 32'hc28891b2;
    11'd1804: sine = 32'hc2881ec6;
    11'd1805: sine = 32'hc287ab87;
    11'd1806: sine = 32'hc28737f3;
    11'd1807: sine = 32'hc286c40c;
    11'd1808: sine = 32'hc2864fd2;
    11'd1809: sine = 32'hc285db46;
    11'd1810: sine = 32'hc2856666;
    11'd1811: sine = 32'hc284f135;
    11'd1812: sine = 32'hc2847bb1;
    11'd1813: sine = 32'hc28405dc;
    11'd1814: sine = 32'hc2838fb5;
    11'd1815: sine = 32'hc283193d;
    11'd1816: sine = 32'hc282a274;
    11'd1817: sine = 32'hc2822b5b;
    11'd1818: sine = 32'hc281b3f1;
    11'd1819: sine = 32'hc2813c37;
    11'd1820: sine = 32'hc280c42e;
    11'd1821: sine = 32'hc2804bd5;
    11'd1822: sine = 32'hc27fa65a;
    11'd1823: sine = 32'hc27eb46c;
    11'd1824: sine = 32'hc27dc1e1;
    11'd1825: sine = 32'hc27cceba;
    11'd1826: sine = 32'hc27bdaf7;
    11'd1827: sine = 32'hc27ae698;
    11'd1828: sine = 32'hc279f19f;
    11'd1829: sine = 32'hc278fc0b;
    11'd1830: sine = 32'hc27805de;
    11'd1831: sine = 32'hc2770f18;
    11'd1832: sine = 32'hc27617b9;
    11'd1833: sine = 32'hc2751fc3;
    11'd1834: sine = 32'hc2742735;
    11'd1835: sine = 32'hc2732e11;
    11'd1836: sine = 32'hc2723457;
    11'd1837: sine = 32'hc2713a07;
    11'd1838: sine = 32'hc2703f23;
    11'd1839: sine = 32'hc26f43aa;
    11'd1840: sine = 32'hc26e479e;
    11'd1841: sine = 32'hc26d4aff;
    11'd1842: sine = 32'hc26c4dcd;
    11'd1843: sine = 32'hc26b500a;
    11'd1844: sine = 32'hc26a51b5;
    11'd1845: sine = 32'hc26952d0;
    11'd1846: sine = 32'hc268535b;
    11'd1847: sine = 32'hc2675357;
    11'd1848: sine = 32'hc26652c4;
    11'd1849: sine = 32'hc26551a3;
    11'd1850: sine = 32'hc2644ff5;
    11'd1851: sine = 32'hc2634dba;
    11'd1852: sine = 32'hc2624af2;
    11'd1853: sine = 32'hc261479f;
    11'd1854: sine = 32'hc26043c1;
    11'd1855: sine = 32'hc25f3f59;
    11'd1856: sine = 32'hc25e3a66;
    11'd1857: sine = 32'hc25d34eb;
    11'd1858: sine = 32'hc25c2ee8;
    11'd1859: sine = 32'hc25b285c;
    11'd1860: sine = 32'hc25a214a;
    11'd1861: sine = 32'hc25919b0;
    11'd1862: sine = 32'hc2581191;
    11'd1863: sine = 32'hc25708ed;
    11'd1864: sine = 32'hc255ffc4;
    11'd1865: sine = 32'hc254f617;
    11'd1866: sine = 32'hc253ebe6;
    11'd1867: sine = 32'hc252e133;
    11'd1868: sine = 32'hc251d5fe;
    11'd1869: sine = 32'hc250ca47;
    11'd1870: sine = 32'hc24fbe10;
    11'd1871: sine = 32'hc24eb158;
    11'd1872: sine = 32'hc24da421;
    11'd1873: sine = 32'hc24c966b;
    11'd1874: sine = 32'hc24b8837;
    11'd1875: sine = 32'hc24a7985;
    11'd1876: sine = 32'hc2496a57;
    11'd1877: sine = 32'hc2485aac;
    11'd1878: sine = 32'hc2474a86;
    11'd1879: sine = 32'hc24639e4;
    11'd1880: sine = 32'hc24528c9;
    11'd1881: sine = 32'hc2441733;
    11'd1882: sine = 32'hc2430525;
    11'd1883: sine = 32'hc241f29f;
    11'd1884: sine = 32'hc240dfa1;
    11'd1885: sine = 32'hc23fcc2b;
    11'd1886: sine = 32'hc23eb840;
    11'd1887: sine = 32'hc23da3df;
    11'd1888: sine = 32'hc23c8f09;
    11'd1889: sine = 32'hc23b79bf;
    11'd1890: sine = 32'hc23a6401;
    11'd1891: sine = 32'hc2394dd0;
    11'd1892: sine = 32'hc238372c;
    11'd1893: sine = 32'hc2372017;
    11'd1894: sine = 32'hc2360892;
    11'd1895: sine = 32'hc234f09b;
    11'd1896: sine = 32'hc233d836;
    11'd1897: sine = 32'hc232bf61;
    11'd1898: sine = 32'hc231a61e;
    11'd1899: sine = 32'hc2308c6d;
    11'd1900: sine = 32'hc22f7250;
    11'd1901: sine = 32'hc22e57c6;
    11'd1902: sine = 32'hc22d3cd1;
    11'd1903: sine = 32'hc22c2171;
    11'd1904: sine = 32'hc22b05a7;
    11'd1905: sine = 32'hc229e973;
    11'd1906: sine = 32'hc228ccd6;
    11'd1907: sine = 32'hc227afd2;
    11'd1908: sine = 32'hc2269265;
    11'd1909: sine = 32'hc2257493;
    11'd1910: sine = 32'hc224565a;
    11'd1911: sine = 32'hc22337bb;
    11'd1912: sine = 32'hc22218b8;
    11'd1913: sine = 32'hc220f951;
    11'd1914: sine = 32'hc21fd987;
    11'd1915: sine = 32'hc21eb95a;
    11'd1916: sine = 32'hc21d98cb;
    11'd1917: sine = 32'hc21c77db;
    11'd1918: sine = 32'hc21b568b;
    11'd1919: sine = 32'hc21a34da;
    11'd1920: sine = 32'hc21912cb;
    11'd1921: sine = 32'hc217f05d;
    11'd1922: sine = 32'hc216cd91;
    11'd1923: sine = 32'hc215aa69;
    11'd1924: sine = 32'hc21486e4;
    11'd1925: sine = 32'hc2136303;
    11'd1926: sine = 32'hc2123ec8;
    11'd1927: sine = 32'hc2111a32;
    11'd1928: sine = 32'hc20ff543;
    11'd1929: sine = 32'hc20ecffb;
    11'd1930: sine = 32'hc20daa5b;
    11'd1931: sine = 32'hc20c8463;
    11'd1932: sine = 32'hc20b5e15;
    11'd1933: sine = 32'hc20a3771;
    11'd1934: sine = 32'hc2091078;
    11'd1935: sine = 32'hc207e92a;
    11'd1936: sine = 32'hc206c188;
    11'd1937: sine = 32'hc2059993;
    11'd1938: sine = 32'hc204714c;
    11'd1939: sine = 32'hc20348b3;
    11'd1940: sine = 32'hc2021fc9;
    11'd1941: sine = 32'hc200f68e;
    11'd1942: sine = 32'hc1ff9a09;
    11'd1943: sine = 32'hc1fd4658;
    11'd1944: sine = 32'hc1faf20a;
    11'd1945: sine = 32'hc1f89d22;
    11'd1946: sine = 32'hc1f647a0;
    11'd1947: sine = 32'hc1f3f187;
    11'd1948: sine = 32'hc1f19ad7;
    11'd1949: sine = 32'hc1ef4392;
    11'd1950: sine = 32'hc1ecebb9;
    11'd1951: sine = 32'hc1ea934e;
    11'd1952: sine = 32'hc1e83a52;
    11'd1953: sine = 32'hc1e5e0c8;
    11'd1954: sine = 32'hc1e386af;
    11'd1955: sine = 32'hc1e12c0a;
    11'd1956: sine = 32'hc1ded0da;
    11'd1957: sine = 32'hc1dc7521;
    11'd1958: sine = 32'hc1da18e0;
    11'd1959: sine = 32'hc1d7bc18;
    11'd1960: sine = 32'hc1d55ecb;
    11'd1961: sine = 32'hc1d300fb;
    11'd1962: sine = 32'hc1d0a2a8;
    11'd1963: sine = 32'hc1ce43d4;
    11'd1964: sine = 32'hc1cbe482;
    11'd1965: sine = 32'hc1c984b2;
    11'd1966: sine = 32'hc1c72465;
    11'd1967: sine = 32'hc1c4c39d;
    11'd1968: sine = 32'hc1c2625c;
    11'd1969: sine = 32'hc1c000a4;
    11'd1970: sine = 32'hc1bd9e74;
    11'd1971: sine = 32'hc1bb3bd0;
    11'd1972: sine = 32'hc1b8d8b9;
    11'd1973: sine = 32'hc1b6752f;
    11'd1974: sine = 32'hc1b41135;
    11'd1975: sine = 32'hc1b1accb;
    11'd1976: sine = 32'hc1af47f4;
    11'd1977: sine = 32'hc1ace2b1;
    11'd1978: sine = 32'hc1aa7d04;
    11'd1979: sine = 32'hc1a816ed;
    11'd1980: sine = 32'hc1a5b06e;
    11'd1981: sine = 32'hc1a34989;
    11'd1982: sine = 32'hc1a0e240;
    11'd1983: sine = 32'hc19e7a93;
    11'd1984: sine = 32'hc19c1285;
    11'd1985: sine = 32'hc199aa16;
    11'd1986: sine = 32'hc1974149;
    11'd1987: sine = 32'hc194d81e;
    11'd1988: sine = 32'hc1926e97;
    11'd1989: sine = 32'hc19004b6;
    11'd1990: sine = 32'hc18d9a7c;
    11'd1991: sine = 32'hc18b2feb;
    11'd1992: sine = 32'hc188c504;
    11'd1993: sine = 32'hc18659c9;
    11'd1994: sine = 32'hc183ee3a;
    11'd1995: sine = 32'hc181825b;
    11'd1996: sine = 32'hc17e2c56;
    11'd1997: sine = 32'hc179535b;
    11'd1998: sine = 32'hc17479c5;
    11'd1999: sine = 32'hc16f9f99;
    11'd2000: sine = 32'hc16ac4d8;
    11'd2001: sine = 32'hc165e987;
    11'd2002: sine = 32'hc1610da8;
    11'd2003: sine = 32'hc15c313f;
    11'd2004: sine = 32'hc157544d;
    11'd2005: sine = 32'hc15276d7;
    11'd2006: sine = 32'hc14d98de;
    11'd2007: sine = 32'hc148ba67;
    11'd2008: sine = 32'hc143db75;
    11'd2009: sine = 32'hc13efc09;
    11'd2010: sine = 32'hc13a1c27;
    11'd2011: sine = 32'hc1353bd3;
    11'd2012: sine = 32'hc1305b0f;
    11'd2013: sine = 32'hc12b79de;
    11'd2014: sine = 32'hc1269844;
    11'd2015: sine = 32'hc121b642;
    11'd2016: sine = 32'hc11cd3dd;
    11'd2017: sine = 32'hc117f117;
    11'd2018: sine = 32'hc1130df4;
    11'd2019: sine = 32'hc10e2a75;
    11'd2020: sine = 32'hc109469f;
    11'd2021: sine = 32'hc1046275;
    11'd2022: sine = 32'hc0fefbf1;
    11'd2023: sine = 32'hc0f5325b;
    11'd2024: sine = 32'hc0eb682d;
    11'd2025: sine = 32'hc0e19d6f;
    11'd2026: sine = 32'hc0d7d225;
    11'd2027: sine = 32'hc0ce0657;
    11'd2028: sine = 32'hc0c43a09;
    11'd2029: sine = 32'hc0ba6d42;
    11'd2030: sine = 32'hc0b0a008;
    11'd2031: sine = 32'hc0a6d261;
    11'd2032: sine = 32'hc09d0453;
    11'd2033: sine = 32'hc09335e5;
    11'd2034: sine = 32'hc089671b;
    11'd2035: sine = 32'hc07f2ffb;
    11'd2036: sine = 32'hc06b9121;
    11'd2037: sine = 32'hc057f1b6;
    11'd2038: sine = 32'hc04451c6;
    11'd2039: sine = 32'hc030b15c;
    11'd2040: sine = 32'hc01d1086;
    11'd2041: sine = 32'hc0096f4f;
    11'd2042: sine = 32'hbfeb9b86;
    11'd2043: sine = 32'hbfc457dd;
    11'd2044: sine = 32'hbf9d13ba;
    11'd2045: sine = 32'hbf6b9e6e;
    11'd2046: sine = 32'hbf1d14d6;
    11'd2047: sine = 32'hbe9d15ba;
  endcase
end
endmodule
